-- Dump 

arch ia32

objects

ioports = io_ports (64k ports)
untyped@e001d000@12 = ut (12 bits)
untyped@e001e000@12 = ut (12 bits)
untyped@e001f000@12 = ut (12 bits)
untyped@e0020000@12 = ut (12 bits)
untyped@e0021000@12 = ut (12 bits)
untyped@e0022000@12 = ut (12 bits)
untyped@e0026000@12 = ut (12 bits)
untyped@e0027000@12 = ut (12 bits)
untyped@e0028000@12 = ut (12 bits)
untyped@e0029000@12 = ut (12 bits)
untyped@e002a000@12 = ut (12 bits)
untyped@e002b000@12 = ut (12 bits)
untyped@e002c000@12 = ut (12 bits)
untyped@e002d000@12 = ut (12 bits)
untyped@e002e000@12 = ut (12 bits)
untyped@e002f000@12 = ut (12 bits)
untyped@e0030000@12 = ut (12 bits)
untyped@e0031000@12 = ut (12 bits)
untyped@e0032000@12 = ut (12 bits)
untyped@e0033000@12 = ut (12 bits)
untyped@e0034000@12 = ut (12 bits)
untyped@e0035000@12 = ut (12 bits)
untyped@e0036000@12 = ut (12 bits)
untyped@e0037000@12 = ut (12 bits)
untyped@e0038000@12 = ut (12 bits)
untyped@e0039000@12 = ut (12 bits)
untyped@e003a000@12 = ut (12 bits)
untyped@e003b000@12 = ut (12 bits)
untyped@e003c000@12 = ut (12 bits)
untyped@e003d000@12 = ut (12 bits)
untyped@e003e000@12 = ut (12 bits)
untyped@e003f000@12 = ut (12 bits)
untyped@e0090000@12 = ut (12 bits)
untyped@e0091000@12 = ut (12 bits)
untyped@e0092000@12 = ut (12 bits)
untyped@e0093000@12 = ut (12 bits)
untyped@e009c000@12 = ut (12 bits)
untyped@e009d000@12 = ut (12 bits)
untyped@e009e000@12 = ut (12 bits)
untyped@e012e000@12 = ut (12 bits)
untyped@e012f000@12 = ut (12 bits)
untyped@e0131000@12 = ut (12 bits)
untyped@e0133000@12 = ut (12 bits)
untyped@e0134000@12 = ut (12 bits)
untyped@e0135000@12 = ut (12 bits)
untyped@e0136000@12 = ut (12 bits)
untyped@e0137000@12 = ut (12 bits)
untyped@e0138000@12 = ut (12 bits)
untyped@e0139000@12 = ut (12 bits)
untyped@e013a000@12 = ut (12 bits)
untyped@e013b000@12 = ut (12 bits)
untyped@e013c000@12 = ut (12 bits)
untyped@e013d000@12 = ut (12 bits)
untyped@e013e000@12 = ut (12 bits)
untyped@e013f000@12 = ut (12 bits)
untyped@e0200000@20 = ut (20 bits)
untyped@e0300000@20 = ut (20 bits)
untyped@e0800000@20 = ut (20 bits)
untyped@e0900000@20 = ut (20 bits)
untyped@e0a00000@20 = ut (20 bits)
untyped@e0b00000@20 = ut (20 bits)
untyped@e0c40000@12 = ut (12 bits)
untyped@e0c41000@12 = ut (12 bits)
untyped@e0c42000@12 = ut (12 bits)
untyped@e0c43000@12 = ut (12 bits)
untyped@e0c44000@12 = ut (12 bits)
untyped@e0c45000@12 = ut (12 bits)
untyped@e0c46000@12 = ut (12 bits)
untyped@e0c47000@12 = ut (12 bits)
untyped@e0c48000@12 = ut (12 bits)
untyped@e0c49000@12 = ut (12 bits)
untyped@e182d000@12 = ut (12 bits)
untyped@e182e000@12 = ut (12 bits)
untyped@e1900000@20 = ut (20 bits)
untyped@e1a00000@20 = ut (20 bits)
untyped@e1b00000@20 = ut (20 bits)
untyped@e1c00000@20 = ut (20 bits)
untyped@e1d00000@20 = ut (20 bits)
untyped@e1e00000@20 = ut (20 bits)
untyped@e1f00000@20 = ut (20 bits)
untyped@e2000000@20 = ut (20 bits)
untyped@e2100000@20 = ut (20 bits)
untyped@e2200000@20 = ut (20 bits)
untyped@e2300000@20 = ut (20 bits)
untyped@e2400000@20 = ut (20 bits)
untyped@e2500000@20 = ut (20 bits)
untyped@e2600000@20 = ut (20 bits)
untyped@e2700000@20 = ut (20 bits)
untyped@e2800000@20 = ut (20 bits)
untyped@e2900000@20 = ut (20 bits)
untyped@e2a00000@20 = ut (20 bits)
untyped@e2b00000@20 = ut (20 bits)
untyped@e2c00000@20 = ut (20 bits)
untyped@e2d00000@20 = ut (20 bits)
untyped@e2e00000@20 = ut (20 bits)
untyped@e2f00000@20 = ut (20 bits)
untyped@e3000000@20 = ut (20 bits)
untyped@e3100000@20 = ut (20 bits)
untyped@e3200000@20 = ut (20 bits)
untyped@e3300000@20 = ut (20 bits)
untyped@e3400000@20 = ut (20 bits)
untyped@e3500000@20 = ut (20 bits)
untyped@e3600000@20 = ut (20 bits)
untyped@e3700000@20 = ut (20 bits)
untyped@e3800000@20 = ut (20 bits)
untyped@e3900000@20 = ut (20 bits)
untyped@e3a00000@20 = ut (20 bits)
untyped@e3b00000@20 = ut (20 bits)
untyped@e3c00000@20 = ut (20 bits)
untyped@e3d00000@20 = ut (20 bits)
untyped@e3e00000@20 = ut (20 bits)
untyped@e3f00000@20 = ut (20 bits)
untyped@e4000000@20 = ut (20 bits)
untyped@e4100000@20 = ut (20 bits)
untyped@e4200000@20 = ut (20 bits)
untyped@e4300000@20 = ut (20 bits)
untyped@e4400000@20 = ut (20 bits)
untyped@e4500000@20 = ut (20 bits)
untyped@e4600000@20 = ut (20 bits)
untyped@e4700000@20 = ut (20 bits)
untyped@e4800000@20 = ut (20 bits)
untyped@e4900000@20 = ut (20 bits)
untyped@e4a00000@20 = ut (20 bits)
untyped@e4b00000@20 = ut (20 bits)
untyped@e4c00000@20 = ut (20 bits)
untyped@e4d00000@20 = ut (20 bits)
untyped@e4e00000@20 = ut (20 bits)
untyped@e4f00000@20 = ut (20 bits)
untyped@e5000000@20 = ut (20 bits)
untyped@e5100000@20 = ut (20 bits)
untyped@e5200000@20 = ut (20 bits)
untyped@e5300000@20 = ut (20 bits)
untyped@e5400000@20 = ut (20 bits)
untyped@e5500000@20 = ut (20 bits)
untyped@e5600000@20 = ut (20 bits)
untyped@e5700000@20 = ut (20 bits)
untyped@e5800000@20 = ut (20 bits)
untyped@e5900000@20 = ut (20 bits)
untyped@e5a00000@20 = ut (20 bits)
untyped@e5b00000@20 = ut (20 bits)
untyped@e5c00000@20 = ut (20 bits)
untyped@e5d00000@20 = ut (20 bits)
untyped@e5e00000@20 = ut (20 bits)
untyped@e5f00000@20 = ut (20 bits)
untyped@e6000000@20 = ut (20 bits)
untyped@e6100000@20 = ut (20 bits)
untyped@e6200000@20 = ut (20 bits)
untyped@e6300000@20 = ut (20 bits)
untyped@e6400000@20 = ut (20 bits)
untyped@e6500000@20 = ut (20 bits)
untyped@e6600000@20 = ut (20 bits)
untyped@e6700000@20 = ut (20 bits)
untyped@e6800000@20 = ut (20 bits)
untyped@e6900000@20 = ut (20 bits)
untyped@e6a00000@20 = ut (20 bits)
untyped@e6b00000@20 = ut (20 bits)
untyped@e6c00000@20 = ut (20 bits)
untyped@e6d00000@20 = ut (20 bits)
untyped@e6e00000@20 = ut (20 bits)
untyped@e6f00000@20 = ut (20 bits)
untyped@e7000000@20 = ut (20 bits)
untyped@e7100000@20 = ut (20 bits)
untyped@e7200000@20 = ut (20 bits)
untyped@e7300000@20 = ut (20 bits)
untyped@e7400000@20 = ut (20 bits)
untyped@e7500000@20 = ut (20 bits)
untyped@e7600000@20 = ut (20 bits)
untyped@e7700000@20 = ut (20 bits)
untyped@e7800000@20 = ut (20 bits)
untyped@e7900000@20 = ut (20 bits)
untyped@e7a00000@20 = ut (20 bits)
untyped@e7b00000@20 = ut (20 bits)
untyped@e7c00000@20 = ut (20 bits)
untyped@e7d00000@20 = ut (20 bits)
untyped@e7e00000@20 = ut (20 bits)
untyped@e7f00000@20 = ut (20 bits)
untyped@e8000000@20 = ut (20 bits)
untyped@e8100000@20 = ut (20 bits)
untyped@e8200000@20 = ut (20 bits)
untyped@e8300000@20 = ut (20 bits)
untyped@e8400000@20 = ut (20 bits)
untyped@e8500000@20 = ut (20 bits)
untyped@e8600000@20 = ut (20 bits)
untyped@e8700000@20 = ut (20 bits)
untyped@e8800000@20 = ut (20 bits)
untyped@e8900000@20 = ut (20 bits)
untyped@e8a00000@20 = ut (20 bits)
untyped@e8b00000@20 = ut (20 bits)
untyped@e8c00000@20 = ut (20 bits)
untyped@e8d00000@20 = ut (20 bits)
untyped@e8e00000@20 = ut (20 bits)
untyped@e8f00000@20 = ut (20 bits)
untyped@e9000000@20 = ut (20 bits)
untyped@e9100000@20 = ut (20 bits)
untyped@e9200000@20 = ut (20 bits)
untyped@e9300000@20 = ut (20 bits)
untyped@e9400000@20 = ut (20 bits)
untyped@e9500000@20 = ut (20 bits)
untyped@e9600000@20 = ut (20 bits)
untyped@e9700000@20 = ut (20 bits)
untyped@e9800000@20 = ut (20 bits)
untyped@e9900000@20 = ut (20 bits)
untyped@e9a00000@20 = ut (20 bits)
untyped@e9b00000@20 = ut (20 bits)
untyped@e9c00000@20 = ut (20 bits)
untyped@e9d00000@20 = ut (20 bits)
untyped@e9e00000@20 = ut (20 bits)
untyped@e9f00000@20 = ut (20 bits)
untyped@ea000000@20 = ut (20 bits)
untyped@ea100000@20 = ut (20 bits)
untyped@ea200000@20 = ut (20 bits)
untyped@ea300000@20 = ut (20 bits)
untyped@ea400000@20 = ut (20 bits)
untyped@ea500000@20 = ut (20 bits)
untyped@ea600000@20 = ut (20 bits)
untyped@ea700000@20 = ut (20 bits)
untyped@ea800000@20 = ut (20 bits)
untyped@ea900000@20 = ut (20 bits)
untyped@eaa00000@20 = ut (20 bits)
untyped@eab00000@20 = ut (20 bits)
untyped@eac00000@20 = ut (20 bits)
untyped@ead00000@20 = ut (20 bits)
untyped@eae00000@20 = ut (20 bits)
untyped@eaf00000@20 = ut (20 bits)
untyped@eb000000@20 = ut (20 bits)
untyped@eb100000@20 = ut (20 bits)
untyped@eb200000@20 = ut (20 bits)
untyped@eb300000@20 = ut (20 bits)
untyped@eb400000@20 = ut (20 bits)
untyped@eb500000@20 = ut (20 bits)
untyped@eb600000@20 = ut (20 bits)
untyped@eb700000@20 = ut (20 bits)
untyped@eb800000@20 = ut (20 bits)
untyped@eb900000@20 = ut (20 bits)
untyped@eba00000@20 = ut (20 bits)
untyped@ebb00000@20 = ut (20 bits)
untyped@ebc00000@20 = ut (20 bits)
untyped@ebd00000@20 = ut (20 bits)
untyped@ebe00000@20 = ut (20 bits)
untyped@ebf00000@20 = ut (20 bits)
untyped@ec000000@20 = ut (20 bits)
untyped@ec100000@20 = ut (20 bits)
untyped@ec200000@20 = ut (20 bits)
untyped@ec300000@20 = ut (20 bits)
untyped@ec400000@20 = ut (20 bits)
untyped@ec500000@20 = ut (20 bits)
untyped@ec600000@20 = ut (20 bits)
untyped@ec700000@20 = ut (20 bits)
untyped@ec800000@20 = ut (20 bits)
untyped@ec900000@20 = ut (20 bits)
untyped@eca00000@20 = ut (20 bits)
untyped@ecb00000@20 = ut (20 bits)
untyped@ecc00000@20 = ut (20 bits)
untyped@ecd00000@20 = ut (20 bits)
untyped@ece00000@20 = ut (20 bits)
untyped@ecf00000@20 = ut (20 bits)
untyped@ed000000@20 = ut (20 bits)
untyped@ed100000@20 = ut (20 bits)
untyped@ed200000@20 = ut (20 bits)
untyped@ed300000@20 = ut (20 bits)
untyped@ed400000@20 = ut (20 bits)
untyped@ed500000@20 = ut (20 bits)
untyped@ed600000@20 = ut (20 bits)
untyped@ed700000@20 = ut (20 bits)
untyped@ed800000@20 = ut (20 bits)
untyped@ed900000@20 = ut (20 bits)
untyped@eda00000@20 = ut (20 bits)
untyped@edb00000@20 = ut (20 bits)
untyped@edc00000@20 = ut (20 bits)
untyped@edd00000@20 = ut (20 bits)
untyped@ede00000@20 = ut (20 bits)
untyped@edf00000@20 = ut (20 bits)
untyped@ee000000@20 = ut (20 bits)
untyped@ee100000@20 = ut (20 bits)
untyped@ee200000@20 = ut (20 bits)
untyped@ee300000@20 = ut (20 bits)
untyped@ee400000@20 = ut (20 bits)
untyped@ee500000@20 = ut (20 bits)
untyped@ee600000@20 = ut (20 bits)
untyped@ee700000@20 = ut (20 bits)
untyped@ee800000@20 = ut (20 bits)
untyped@ee900000@20 = ut (20 bits)
untyped@eea00000@20 = ut (20 bits)
untyped@eeb00000@20 = ut (20 bits)
untyped@eec00000@20 = ut (20 bits)
untyped@eed00000@20 = ut (20 bits)
untyped@eee00000@20 = ut (20 bits)
untyped@eef00000@20 = ut (20 bits)
untyped@ef000000@20 = ut (20 bits)
untyped@ef100000@20 = ut (20 bits)
untyped@ef200000@20 = ut (20 bits)
untyped@f7300000@20 = ut (20 bits)
untyped@f7400000@20 = ut (20 bits)
untyped@f7500000@20 = ut (20 bits)
untyped@f7600000@20 = ut (20 bits)
untyped@f7700000@20 = ut (20 bits)
untyped@f7800000@20 = ut (20 bits)
untyped@f7900000@20 = ut (20 bits)
untyped@f7a00000@20 = ut (20 bits)
untyped@f7b00000@20 = ut (20 bits)
untyped@f7c00000@20 = ut (20 bits)
untyped@f7d00000@20 = ut (20 bits)
untyped@f7e00000@20 = ut (20 bits)
untyped@f7f00000@20 = ut (20 bits)
untyped@f8000000@20 = ut (20 bits)
untyped@f8100000@20 = ut (20 bits)
untyped@f8200000@20 = ut (20 bits)
untyped@f8300000@20 = ut (20 bits)
untyped@f8400000@20 = ut (20 bits)
untyped@f8500000@20 = ut (20 bits)
untyped@f8600000@20 = ut (20 bits)
untyped@f8700000@20 = ut (20 bits)
untyped@f8800000@20 = ut (20 bits)
untyped@f8900000@20 = ut (20 bits)
untyped@f8a00000@20 = ut (20 bits)
untyped@f8b00000@20 = ut (20 bits)
untyped@f8c00000@20 = ut (20 bits)
untyped@f8d00000@20 = ut (20 bits)
untyped@f8e00000@20 = ut (20 bits)
untyped@f8f00000@20 = ut (20 bits)
untyped@f9000000@20 = ut (20 bits)
untyped@f9100000@20 = ut (20 bits)
untyped@f9200000@20 = ut (20 bits)
untyped@f9300000@20 = ut (20 bits)
untyped@f9400000@20 = ut (20 bits)
untyped@f9500000@20 = ut (20 bits)
untyped@f9600000@20 = ut (20 bits)
untyped@f9700000@20 = ut (20 bits)
untyped@f9e00000@20 = ut (20 bits)
untyped@f9f00000@20 = ut (20 bits)
untyped@fa000000@20 = ut (20 bits)
untyped@fa100000@20 = ut (20 bits)
untyped@fa200000@20 = ut (20 bits)
untyped@fa300000@20 = ut (20 bits)
untyped@fa400000@20 = ut (20 bits)
untyped@fa500000@20 = ut (20 bits)
untyped@fa600000@20 = ut (20 bits)
untyped@fa700000@20 = ut (20 bits)
untyped@fa800000@20 = ut (20 bits)
untyped@fa900000@20 = ut (20 bits)
untyped@faa00000@20 = ut (20 bits)
untyped@fab00000@20 = ut (20 bits)
untyped@fac00000@20 = ut (20 bits)
untyped@fad00000@20 = ut (20 bits)
untyped@fae00000@20 = ut (20 bits)
untyped@faf00000@20 = ut (20 bits)
untyped@fb000000@20 = ut (20 bits)
untyped@fb100000@20 = ut (20 bits)
untyped@fb200000@20 = ut (20 bits)
untyped@fb300000@20 = ut (20 bits)
untyped@fb400000@20 = ut (20 bits)
untyped@fb500000@20 = ut (20 bits)
untyped@fb600000@20 = ut (20 bits)
untyped@fb700000@20 = ut (20 bits)
untyped@fb800000@20 = ut (20 bits)
untyped@fb900000@20 = ut (20 bits)
untyped@fba00000@20 = ut (20 bits)
untyped@fbb00000@20 = ut (20 bits)
untyped@fbc00000@20 = ut (20 bits)
untyped@fbd00000@20 = ut (20 bits)
untyped@fbe00000@20 = ut (20 bits)
untyped@fbf00000@20 = ut (20 bits)
untyped@fc000000@20 = ut (20 bits)
untyped@fc100000@20 = ut (20 bits)
untyped@fc200000@20 = ut (20 bits)
untyped@fc300000@20 = ut (20 bits)
untyped@fc400000@20 = ut (20 bits)
untyped@fc500000@20 = ut (20 bits)
untyped@fc600000@20 = ut (20 bits)
untyped@fc700000@20 = ut (20 bits)
untyped@fc800000@20 = ut (20 bits)
untyped@fc900000@20 = ut (20 bits)
untyped@fca00000@20 = ut (20 bits)
untyped@fcb00000@20 = ut (20 bits)
untyped@fcc00000@20 = ut (20 bits)
untyped@fcd00000@20 = ut (20 bits)
untyped@fce00000@20 = ut (20 bits)
untyped@fcf00000@20 = ut (20 bits)
untyped@fd000000@20 = ut (20 bits)
untyped@fd100000@20 = ut (20 bits)
untyped@fd200000@20 = ut (20 bits)
untyped@fd300000@20 = ut (20 bits)
untyped@fd400000@20 = ut (20 bits)
untyped@fd500000@20 = ut (20 bits)
untyped@fd600000@20 = ut (20 bits)
untyped@fd700000@20 = ut (20 bits)
untyped@fd800000@20 = ut (20 bits)
untyped@fd900000@20 = ut (20 bits)
untyped@fda00000@20 = ut (20 bits)
untyped@fdb00000@20 = ut (20 bits)
untyped@fdc00000@20 = ut (20 bits)
untyped@fdd00000@20 = ut (20 bits)
untyped@fde00000@20 = ut (20 bits)
untyped@fdf00000@20 = ut (20 bits)
untyped@fe000000@20 = ut (20 bits)
untyped@fe100000@20 = ut (20 bits)
untyped@fe200000@20 = ut (20 bits)
untyped@fe300000@20 = ut (20 bits)
untyped@fe400000@20 = ut (20 bits)
untyped@fe500000@20 = ut (20 bits)
untyped@fe600000@20 = ut (20 bits)
untyped@fe700000@20 = ut (20 bits)
untyped@fe800000@20 = ut (20 bits)
untyped@fe900000@20 = ut (20 bits)
untyped@fea00000@20 = ut (20 bits)
untyped@feb00000@20 = ut (20 bits)
untyped@fec00000@20 = ut (20 bits)
untyped@fed00000@20 = ut (20 bits)
untyped@fee00000@20 = ut (20 bits)
untyped@fef00000@20 = ut (20 bits)
untyped@ff000000@20 = ut (20 bits)
untyped@ff100000@20 = ut (20 bits)
untyped@ff200000@20 = ut (20 bits)
untyped@ff300000@20 = ut (20 bits)
untyped@ff400000@20 = ut (20 bits)
untyped@ff500000@20 = ut (20 bits)
untyped@ff600000@20 = ut (20 bits)
untyped@ff700000@20 = ut (20 bits)
untyped@ff800000@20 = ut (20 bits)
untyped@ff900000@20 = ut (20 bits)
untyped@ffa00000@20 = ut (20 bits)
untyped@ffb00000@20 = ut (20 bits)
untyped@ffc00000@20 = ut (20 bits)
untyped@ffd00000@20 = ut (20 bits)
ep@e001cff0 = ep
aep@fffeffd0 = aep
aep@fffeffe0 = aep
cnode@f6bc8000 = cnode(10 bits) 
cnode@f6bcc000 = cnode(10 bits) 
cnode@f6bf0000 = cnode(10 bits) 
cnode@f6bf4000 = cnode(10 bits) 
tcb@fffee500 = tcb
tcb@fffee900 = tcb
tcb@fffeed00 = tcb
frame@d0180000 = frame(4k)
frame@d0181000 = frame(4k)
frame@d0182000 = frame(4k)
frame@d0183000 = frame(4k)
frame@d0184000 = frame(4k)
frame@d0185000 = frame(4k)
frame@d0186000 = frame(4k)
frame@d0187000 = frame(4k)
frame@d0188000 = frame(4k)
frame@d0189000 = frame(4k)
frame@d018a000 = frame(4k)
frame@d018b000 = frame(4k)
frame@d018c000 = frame(4k)
frame@d018d000 = frame(4k)
frame@d018e000 = frame(4k)
frame@d018f000 = frame(4k)
frame@d0190000 = frame(4k)
frame@d0191000 = frame(4k)
frame@d0192000 = frame(4k)
frame@d0193000 = frame(4k)
frame@d0194000 = frame(4k)
frame@d0195000 = frame(4k)
frame@d0196000 = frame(4k)
frame@d0197000 = frame(4k)
frame@d0198000 = frame(4k)
frame@d0199000 = frame(4k)
frame@d019a000 = frame(4k)
frame@d019b000 = frame(4k)
frame@d019c000 = frame(4k)
frame@d019d000 = frame(4k)
frame@d019e000 = frame(4k)
frame@d019f000 = frame(4k)
frame@d01a5000 = frame(4k)
frame@d0200000 = frame(4k)
frame@d0201000 = frame(4k)
frame@d0202000 = frame(4k)
frame@d0203000 = frame(4k)
frame@d0204000 = frame(4k)
frame@d0205000 = frame(4k)
frame@d0206000 = frame(4k)
frame@d0207000 = frame(4k)
frame@d0208000 = frame(4k)
frame@d0209000 = frame(4k)
frame@d020a000 = frame(4k)
frame@d020b000 = frame(4k)
frame@d020c000 = frame(4k)
frame@d020d000 = frame(4k)
frame@d020e000 = frame(4k)
frame@d020f000 = frame(4k)
frame@d0210000 = frame(4k)
frame@d0211000 = frame(4k)
frame@d0212000 = frame(4k)
frame@d0213000 = frame(4k)
frame@d0214000 = frame(4k)
frame@d0215000 = frame(4k)
frame@d0216000 = frame(4k)
frame@d0217000 = frame(4k)
frame@d0218000 = frame(4k)
frame@d0219000 = frame(4k)
frame@d021a000 = frame(4k)
frame@d021b000 = frame(4k)
frame@d021c000 = frame(4k)
frame@d021d000 = frame(4k)
frame@d021e000 = frame(4k)
frame@d021f000 = frame(4k)
frame@d0220000 = frame(4k)
frame@d0221000 = frame(4k)
frame@d0222000 = frame(4k)
frame@d0223000 = frame(4k)
frame@d0224000 = frame(4k)
frame@d0225000 = frame(4k)
frame@d0226000 = frame(4k)
frame@d0227000 = frame(4k)
frame@d0228000 = frame(4k)
frame@d0229000 = frame(4k)
frame@d022a000 = frame(4k)
frame@d022b000 = frame(4k)
frame@d022c000 = frame(4k)
frame@d022d000 = frame(4k)
frame@d022e000 = frame(4k)
frame@d022f000 = frame(4k)
frame@d0230000 = frame(4k)
frame@d0231000 = frame(4k)
frame@d0232000 = frame(4k)
frame@d0233000 = frame(4k)
frame@d0234000 = frame(4k)
frame@d0235000 = frame(4k)
frame@d0236000 = frame(4k)
frame@d0237000 = frame(4k)
frame@d0238000 = frame(4k)
frame@d0239000 = frame(4k)
frame@d023a000 = frame(4k)
frame@d023b000 = frame(4k)
frame@d023c000 = frame(4k)
frame@d023d000 = frame(4k)
frame@d023e000 = frame(4k)
frame@d023f000 = frame(4k)
frame@d0240000 = frame(4k)
frame@d0241000 = frame(4k)
frame@d0242000 = frame(4k)
frame@d0243000 = frame(4k)
frame@d0244000 = frame(4k)
frame@d0245000 = frame(4k)
frame@d0246000 = frame(4k)
frame@d0247000 = frame(4k)
frame@d0248000 = frame(4k)
frame@d0249000 = frame(4k)
frame@d024a000 = frame(4k)
frame@d024b000 = frame(4k)
frame@d024c000 = frame(4k)
frame@d024d000 = frame(4k)
frame@d024e000 = frame(4k)
frame@d024f000 = frame(4k)
frame@d0250000 = frame(4k)
frame@d0251000 = frame(4k)
frame@d0252000 = frame(4k)
frame@d0253000 = frame(4k)
frame@d0254000 = frame(4k)
frame@d0255000 = frame(4k)
frame@d0256000 = frame(4k)
frame@d0257000 = frame(4k)
frame@d0258000 = frame(4k)
frame@d0259000 = frame(4k)
frame@d025a000 = frame(4k)
frame@d025b000 = frame(4k)
frame@d025c000 = frame(4k)
frame@d025d000 = frame(4k)
frame@d025e000 = frame(4k)
frame@d025f000 = frame(4k)
frame@d0260000 = frame(4k)
frame@d0261000 = frame(4k)
frame@d0262000 = frame(4k)
frame@d0263000 = frame(4k)
frame@d0264000 = frame(4k)
frame@d0265000 = frame(4k)
frame@d0266000 = frame(4k)
frame@d0267000 = frame(4k)
frame@d0268000 = frame(4k)
frame@d0269000 = frame(4k)
frame@d026a000 = frame(4k)
frame@d026b000 = frame(4k)
frame@d026c000 = frame(4k)
frame@d026d000 = frame(4k)
frame@d026e000 = frame(4k)
frame@d026f000 = frame(4k)
frame@d0270000 = frame(4k)
frame@d0271000 = frame(4k)
frame@d0272000 = frame(4k)
frame@d0273000 = frame(4k)
frame@d0274000 = frame(4k)
frame@d0275000 = frame(4k)
frame@d0276000 = frame(4k)
frame@d0277000 = frame(4k)
frame@d0278000 = frame(4k)
frame@d0279000 = frame(4k)
frame@d027a000 = frame(4k)
frame@d027b000 = frame(4k)
frame@d027c000 = frame(4k)
frame@d027d000 = frame(4k)
frame@d027e000 = frame(4k)
frame@d027f000 = frame(4k)
frame@d0300000 = frame(4k)
frame@d0301000 = frame(4k)
frame@d0302000 = frame(4k)
frame@d0303000 = frame(4k)
frame@f6c80000 = frame(4k)
frame@f6c81000 = frame(4k)
frame@f6c82000 = frame(4k)
frame@f6c83000 = frame(4k)
frame@f6c84000 = frame(4k)
frame@f6c85000 = frame(4k)
frame@f6c86000 = frame(4k)
frame@f6c87000 = frame(4k)
frame@f6c88000 = frame(4k)
frame@f6c89000 = frame(4k)
frame@f6c8a000 = frame(4k)
frame@f6c8b000 = frame(4k)
frame@f6c8c000 = frame(4k)
frame@f6c8d000 = frame(4k)
frame@f6c8e000 = frame(4k)
frame@f6c8f000 = frame(4k)
frame@f6c90000 = frame(4k)
frame@f6c91000 = frame(4k)
frame@f6c92000 = frame(4k)
frame@f6c93000 = frame(4k)
frame@f6c94000 = frame(4k)
frame@f6c95000 = frame(4k)
frame@f6c96000 = frame(4k)
frame@f6c97000 = frame(4k)
frame@f6c98000 = frame(4k)
frame@f6c99000 = frame(4k)
frame@f6c9a000 = frame(4k)
frame@f6c9b000 = frame(4k)
frame@f6c9c000 = frame(4k)
frame@f6c9d000 = frame(4k)
frame@f6c9e000 = frame(4k)
frame@f6c9f000 = frame(4k)
frame@f6ca0000 = frame(4k)
frame@f6ca1000 = frame(4k)
frame@f6ca2000 = frame(4k)
frame@f6ca3000 = frame(4k)
frame@f6ca4000 = frame(4k)
frame@f6ca5000 = frame(4k)
frame@f6ca6000 = frame(4k)
frame@f6ca7000 = frame(4k)
frame@f6ca8000 = frame(4k)
frame@f6ca9000 = frame(4k)
frame@f6caa000 = frame(4k)
frame@f6cab000 = frame(4k)
frame@f6cac000 = frame(4k)
frame@f6cad000 = frame(4k)
frame@f6cae000 = frame(4k)
frame@f6caf000 = frame(4k)
frame@f6cb0000 = frame(4k)
frame@f6cb1000 = frame(4k)
frame@f6cb2000 = frame(4k)
frame@f6cb3000 = frame(4k)
frame@f6cb4000 = frame(4k)
frame@f6cb5000 = frame(4k)
frame@f6cb6000 = frame(4k)
frame@f6cb7000 = frame(4k)
frame@f6cb8000 = frame(4k)
frame@f6cb9000 = frame(4k)
frame@f6cba000 = frame(4k)
frame@f6cbb000 = frame(4k)
frame@f6cbc000 = frame(4k)
frame@f6cbd000 = frame(4k)
frame@f6cbe000 = frame(4k)
frame@f6cbf000 = frame(4k)
frame@f6cc0000 = frame(4k)
frame@f6cc1000 = frame(4k)
frame@f6cc2000 = frame(4k)
frame@f6cc3000 = frame(4k)
frame@f6cc4000 = frame(4k)
frame@f6cc5000 = frame(4k)
frame@f6cc6000 = frame(4k)
frame@f6cc7000 = frame(4k)
frame@f6cc8000 = frame(4k)
frame@f6cc9000 = frame(4k)
frame@f6cca000 = frame(4k)
frame@f6ccb000 = frame(4k)
frame@f6ccc000 = frame(4k)
frame@f6ccd000 = frame(4k)
frame@f6cce000 = frame(4k)
frame@f6ccf000 = frame(4k)
frame@f6cd0000 = frame(4k)
frame@f6cd1000 = frame(4k)
frame@f6cd2000 = frame(4k)
frame@f6cd3000 = frame(4k)
frame@f6cd4000 = frame(4k)
frame@f6cd5000 = frame(4k)
frame@f6cd6000 = frame(4k)
frame@f6cd7000 = frame(4k)
frame@f6cd8000 = frame(4k)
frame@f6cd9000 = frame(4k)
frame@f6cda000 = frame(4k)
frame@f6cdb000 = frame(4k)
frame@f6cdc000 = frame(4k)
frame@f6cdd000 = frame(4k)
frame@f6cde000 = frame(4k)
frame@f6cdf000 = frame(4k)
frame@f6ce0000 = frame(4k)
frame@f6ce1000 = frame(4k)
frame@f6ce2000 = frame(4k)
frame@f6ce3000 = frame(4k)
frame@f6ce4000 = frame(4k)
frame@f6ce5000 = frame(4k)
frame@f6ce6000 = frame(4k)
frame@f6ce7000 = frame(4k)
frame@f6ce8000 = frame(4k)
frame@f6ce9000 = frame(4k)
frame@f6cea000 = frame(4k)
frame@f6ceb000 = frame(4k)
frame@f6cec000 = frame(4k)
frame@f6ced000 = frame(4k)
frame@f6cee000 = frame(4k)
frame@f6cef000 = frame(4k)
frame@f6cf0000 = frame(4k)
frame@f6cf1000 = frame(4k)
frame@f6cf2000 = frame(4k)
frame@f6cf3000 = frame(4k)
frame@f6cf4000 = frame(4k)
frame@f6cf5000 = frame(4k)
frame@f6cf6000 = frame(4k)
frame@f6cf7000 = frame(4k)
frame@f6cf8000 = frame(4k)
frame@f6cf9000 = frame(4k)
frame@f6cfa000 = frame(4k)
frame@f6cfb000 = frame(4k)
frame@f6cfc000 = frame(4k)
frame@f6cfd000 = frame(4k)
frame@f6cfe000 = frame(4k)
frame@f6cff000 = frame(4k)
frame@f6d00000 = frame(4k)
frame@f6d01000 = frame(4k)
frame@f6d02000 = frame(4k)
frame@f6d03000 = frame(4k)
frame@f6d04000 = frame(4k)
frame@f6d05000 = frame(4k)
frame@f6d06000 = frame(4k)
frame@f6d07000 = frame(4k)
frame@f6d08000 = frame(4k)
frame@f6d09000 = frame(4k)
frame@f6d0a000 = frame(4k)
frame@f6d0b000 = frame(4k)
frame@f6d0c000 = frame(4k)
frame@f6d0d000 = frame(4k)
frame@f6d0e000 = frame(4k)
frame@f6d0f000 = frame(4k)
frame@f6d10000 = frame(4k)
frame@f6d11000 = frame(4k)
frame@f6d12000 = frame(4k)
frame@f6d13000 = frame(4k)
frame@f6d14000 = frame(4k)
frame@f6d15000 = frame(4k)
frame@f6d16000 = frame(4k)
frame@f6d17000 = frame(4k)
frame@f6d18000 = frame(4k)
frame@f6d19000 = frame(4k)
frame@f6d1a000 = frame(4k)
frame@f6d1b000 = frame(4k)
frame@f6d1c000 = frame(4k)
frame@f6d1d000 = frame(4k)
frame@f6d1e000 = frame(4k)
frame@f6d1f000 = frame(4k)
frame@f6d20000 = frame(4k)
frame@f6d21000 = frame(4k)
frame@f6d22000 = frame(4k)
frame@f6d23000 = frame(4k)
frame@f6d24000 = frame(4k)
frame@f6d25000 = frame(4k)
frame@f6d26000 = frame(4k)
frame@f6d27000 = frame(4k)
frame@f6d28000 = frame(4k)
frame@f6d29000 = frame(4k)
frame@f6d2a000 = frame(4k)
frame@f6d2b000 = frame(4k)
frame@f6d2c000 = frame(4k)
frame@f6d2d000 = frame(4k)
frame@f6d2e000 = frame(4k)
frame@f6d2f000 = frame(4k)
frame@f6d30000 = frame(4k)
frame@f6d31000 = frame(4k)
frame@f6d32000 = frame(4k)
frame@f6d33000 = frame(4k)
frame@f6d34000 = frame(4k)
frame@f6d35000 = frame(4k)
frame@f6d36000 = frame(4k)
frame@f6d37000 = frame(4k)
frame@f6d38000 = frame(4k)
frame@f6d39000 = frame(4k)
frame@f6d3a000 = frame(4k)
frame@f6d3b000 = frame(4k)
frame@f6d3c000 = frame(4k)
frame@f6d3d000 = frame(4k)
frame@f6d3e000 = frame(4k)
frame@f6d3f000 = frame(4k)
frame@f6d40000 = frame(4k)
frame@f6d41000 = frame(4k)
frame@f6d42000 = frame(4k)
frame@f6d43000 = frame(4k)
frame@f6d44000 = frame(4k)
frame@f6d45000 = frame(4k)
frame@f6d46000 = frame(4k)
frame@f6d47000 = frame(4k)
frame@f6d48000 = frame(4k)
frame@f6d49000 = frame(4k)
frame@f6d4a000 = frame(4k)
frame@f6d4b000 = frame(4k)
frame@f6d4c000 = frame(4k)
frame@f6d4d000 = frame(4k)
frame@f6d4e000 = frame(4k)
frame@f6d4f000 = frame(4k)
frame@f6d50000 = frame(4k)
frame@f6d51000 = frame(4k)
frame@f6d52000 = frame(4k)
frame@f6d53000 = frame(4k)
frame@f6d54000 = frame(4k)
frame@f6d55000 = frame(4k)
frame@f6d56000 = frame(4k)
frame@f6d57000 = frame(4k)
frame@f6d58000 = frame(4k)
frame@f6d59000 = frame(4k)
frame@f6d5a000 = frame(4k)
frame@f6d5b000 = frame(4k)
frame@f6d5c000 = frame(4k)
frame@f6d5d000 = frame(4k)
frame@f6d5e000 = frame(4k)
frame@f6d5f000 = frame(4k)
frame@f6d60000 = frame(4k)
frame@f6d61000 = frame(4k)
frame@f6d62000 = frame(4k)
frame@f6d63000 = frame(4k)
frame@f6d64000 = frame(4k)
frame@f6d65000 = frame(4k)
frame@f6d66000 = frame(4k)
frame@f6d67000 = frame(4k)
frame@f6d68000 = frame(4k)
frame@f6d69000 = frame(4k)
frame@f6d6a000 = frame(4k)
frame@f6d6b000 = frame(4k)
frame@f6d6c000 = frame(4k)
frame@f6d6d000 = frame(4k)
frame@f6d6e000 = frame(4k)
frame@f6d6f000 = frame(4k)
frame@f6d70000 = frame(4k)
frame@f6d71000 = frame(4k)
frame@f6d72000 = frame(4k)
frame@f6d73000 = frame(4k)
frame@f6d74000 = frame(4k)
frame@f6d75000 = frame(4k)
frame@f6d76000 = frame(4k)
frame@f6d77000 = frame(4k)
frame@f6d78000 = frame(4k)
frame@f6d79000 = frame(4k)
frame@f6d7a000 = frame(4k)
frame@f6d7b000 = frame(4k)
frame@f6d7c000 = frame(4k)
frame@f6d7d000 = frame(4k)
frame@f6d7e000 = frame(4k)
frame@f6d7f000 = frame(4k)
frame@f6e00000 = frame(4k)
frame@f6e01000 = frame(4k)
frame@f6e02000 = frame(4k)
frame@f6e03000 = frame(4k)
frame@f6e04000 = frame(4k)
frame@f6e05000 = frame(4k)
frame@f6e06000 = frame(4k)
frame@f6e07000 = frame(4k)
frame@f6e08000 = frame(4k)
frame@f6e09000 = frame(4k)
frame@f6e0a000 = frame(4k)
frame@f6e0b000 = frame(4k)
frame@f6e0c000 = frame(4k)
frame@f6e0d000 = frame(4k)
frame@f6e0e000 = frame(4k)
frame@f6e0f000 = frame(4k)
frame@f6e10000 = frame(4k)
frame@f6e11000 = frame(4k)
frame@f6e12000 = frame(4k)
frame@f6e13000 = frame(4k)
frame@f6e14000 = frame(4k)
frame@f6e15000 = frame(4k)
frame@f6e16000 = frame(4k)
frame@f6e17000 = frame(4k)
frame@f6e18000 = frame(4k)
frame@f6e19000 = frame(4k)
frame@f6e1a000 = frame(4k)
frame@f6e1b000 = frame(4k)
frame@f6e1c000 = frame(4k)
frame@f6e1d000 = frame(4k)
frame@f6e1e000 = frame(4k)
frame@f6e1f000 = frame(4k)
frame@f6e20000 = frame(4k)
frame@f6e21000 = frame(4k)
frame@f6e22000 = frame(4k)
frame@f6e23000 = frame(4k)
frame@f6e24000 = frame(4k)
frame@f6e25000 = frame(4k)
frame@f6e26000 = frame(4k)
frame@f6e27000 = frame(4k)
frame@f6e28000 = frame(4k)
frame@f6e29000 = frame(4k)
frame@f6e2a000 = frame(4k)
frame@f6e2b000 = frame(4k)
frame@f6e2c000 = frame(4k)
frame@f6e2d000 = frame(4k)
frame@f6e2e000 = frame(4k)
frame@f6e2f000 = frame(4k)
frame@f6e30000 = frame(4k)
frame@f6e31000 = frame(4k)
frame@f6e32000 = frame(4k)
frame@f6e33000 = frame(4k)
frame@f6e34000 = frame(4k)
frame@f6e35000 = frame(4k)
frame@f6e36000 = frame(4k)
frame@f6e37000 = frame(4k)
frame@f6e38000 = frame(4k)
frame@f6e39000 = frame(4k)
frame@f6e3a000 = frame(4k)
frame@f6e3b000 = frame(4k)
frame@f6e3c000 = frame(4k)
frame@f6e3d000 = frame(4k)
frame@f6e3e000 = frame(4k)
frame@f6e3f000 = frame(4k)
frame@f6e40000 = frame(4k)
frame@f6e41000 = frame(4k)
frame@f6e42000 = frame(4k)
frame@f6e43000 = frame(4k)
frame@f6e44000 = frame(4k)
frame@f6e45000 = frame(4k)
frame@f6e46000 = frame(4k)
frame@f6e47000 = frame(4k)
frame@f6e48000 = frame(4k)
frame@f6e49000 = frame(4k)
frame@f6e4a000 = frame(4k)
frame@f6e4b000 = frame(4k)
frame@f6e4c000 = frame(4k)
frame@f6e4d000 = frame(4k)
frame@f6e4e000 = frame(4k)
frame@f6e4f000 = frame(4k)
frame@f6e50000 = frame(4k)
frame@f6e51000 = frame(4k)
frame@f6e52000 = frame(4k)
frame@f6e53000 = frame(4k)
frame@f6e54000 = frame(4k)
frame@f6e55000 = frame(4k)
frame@f6e56000 = frame(4k)
frame@f6e57000 = frame(4k)
frame@f6e58000 = frame(4k)
frame@f6e59000 = frame(4k)
frame@f6e5a000 = frame(4k)
frame@f6e5b000 = frame(4k)
frame@f6e5c000 = frame(4k)
frame@f6e5d000 = frame(4k)
frame@f6e5e000 = frame(4k)
frame@f6e5f000 = frame(4k)
frame@f6e60000 = frame(4k)
frame@f6e61000 = frame(4k)
frame@f6e62000 = frame(4k)
frame@f6e63000 = frame(4k)
frame@f6e64000 = frame(4k)
frame@f6e65000 = frame(4k)
frame@f6e66000 = frame(4k)
frame@f6e67000 = frame(4k)
frame@f6e68000 = frame(4k)
frame@f6e69000 = frame(4k)
frame@f6e6a000 = frame(4k)
frame@f6e6b000 = frame(4k)
frame@f6e6c000 = frame(4k)
frame@f6e6d000 = frame(4k)
frame@f6e6e000 = frame(4k)
frame@f6e6f000 = frame(4k)
frame@f6e70000 = frame(4k)
frame@f6e71000 = frame(4k)
frame@f6e72000 = frame(4k)
frame@f6e73000 = frame(4k)
frame@f6e74000 = frame(4k)
frame@f6e75000 = frame(4k)
frame@f6e76000 = frame(4k)
frame@f6e77000 = frame(4k)
frame@f6e78000 = frame(4k)
frame@f6e79000 = frame(4k)
frame@f6e7a000 = frame(4k)
frame@f6e7b000 = frame(4k)
frame@f6e7c000 = frame(4k)
frame@f6e7d000 = frame(4k)
frame@f6e7e000 = frame(4k)
frame@f6e7f000 = frame(4k)
frame@f6e80000 = frame(4k)
frame@f6e81000 = frame(4k)
frame@f6e82000 = frame(4k)
frame@f6e83000 = frame(4k)
frame@f6e84000 = frame(4k)
frame@f6e85000 = frame(4k)
frame@f6e86000 = frame(4k)
frame@f6e87000 = frame(4k)
frame@f6e88000 = frame(4k)
frame@f6e89000 = frame(4k)
frame@f6e8a000 = frame(4k)
frame@f6e8b000 = frame(4k)
frame@f6e8c000 = frame(4k)
frame@f6e8d000 = frame(4k)
frame@f6e8e000 = frame(4k)
frame@f6e8f000 = frame(4k)
frame@f6e90000 = frame(4k)
frame@f6e91000 = frame(4k)
frame@f6e92000 = frame(4k)
frame@f6e93000 = frame(4k)
frame@f6e94000 = frame(4k)
frame@f6e95000 = frame(4k)
frame@f6e96000 = frame(4k)
frame@f6e97000 = frame(4k)
frame@f6e98000 = frame(4k)
frame@f6e99000 = frame(4k)
frame@f6e9a000 = frame(4k)
frame@f6e9b000 = frame(4k)
frame@f6e9c000 = frame(4k)
frame@f6e9d000 = frame(4k)
frame@f6e9e000 = frame(4k)
frame@f6e9f000 = frame(4k)
frame@f6ea0000 = frame(4k)
frame@f6ea1000 = frame(4k)
frame@f6ea2000 = frame(4k)
frame@f6ea3000 = frame(4k)
frame@f6ea4000 = frame(4k)
frame@f6ea5000 = frame(4k)
frame@f6ea6000 = frame(4k)
frame@f6ea7000 = frame(4k)
frame@f6ea8000 = frame(4k)
frame@f6ea9000 = frame(4k)
frame@f6eaa000 = frame(4k)
frame@f6eab000 = frame(4k)
frame@f6eac000 = frame(4k)
frame@f6ead000 = frame(4k)
frame@f6eae000 = frame(4k)
frame@f6eaf000 = frame(4k)
frame@f6eb0000 = frame(4k)
frame@f6eb1000 = frame(4k)
frame@f6eb2000 = frame(4k)
frame@f6eb3000 = frame(4k)
frame@f6eb4000 = frame(4k)
frame@f6eb5000 = frame(4k)
frame@f6eb6000 = frame(4k)
frame@f6eb7000 = frame(4k)
frame@f6eb8000 = frame(4k)
frame@f6eb9000 = frame(4k)
frame@f6eba000 = frame(4k)
frame@f6ebb000 = frame(4k)
frame@f6ebc000 = frame(4k)
frame@f6ebd000 = frame(4k)
frame@f6ebe000 = frame(4k)
frame@f6ebf000 = frame(4k)
frame@f6ec0000 = frame(4k)
frame@f6ec1000 = frame(4k)
frame@f6ec2000 = frame(4k)
frame@f6ec3000 = frame(4k)
frame@f6ec4000 = frame(4k)
frame@f6ec5000 = frame(4k)
frame@f6ec6000 = frame(4k)
frame@f6ec7000 = frame(4k)
frame@f6ec8000 = frame(4k)
frame@f6ec9000 = frame(4k)
frame@f6eca000 = frame(4k)
frame@f6ecb000 = frame(4k)
frame@f6ecc000 = frame(4k)
frame@f6ecd000 = frame(4k)
frame@f6ece000 = frame(4k)
frame@f6ecf000 = frame(4k)
frame@f6ed0000 = frame(4k)
frame@f6ed1000 = frame(4k)
frame@f6ed2000 = frame(4k)
frame@f6ed3000 = frame(4k)
frame@f6ed4000 = frame(4k)
frame@f6ed5000 = frame(4k)
frame@f6ed6000 = frame(4k)
frame@f6ed7000 = frame(4k)
frame@f6ed8000 = frame(4k)
frame@f6ed9000 = frame(4k)
frame@f6eda000 = frame(4k)
frame@f6edb000 = frame(4k)
frame@f6edc000 = frame(4k)
frame@f6edd000 = frame(4k)
frame@f6ede000 = frame(4k)
frame@f6edf000 = frame(4k)
frame@f6ee0000 = frame(4k)
frame@f6ee1000 = frame(4k)
frame@f6ee2000 = frame(4k)
frame@f6ee3000 = frame(4k)
frame@f6ee4000 = frame(4k)
frame@f6ee5000 = frame(4k)
frame@f6ee6000 = frame(4k)
frame@f6ee7000 = frame(4k)
frame@f6ee8000 = frame(4k)
frame@f6ee9000 = frame(4k)
frame@f6eea000 = frame(4k)
frame@f6eeb000 = frame(4k)
frame@f6eec000 = frame(4k)
frame@f6eed000 = frame(4k)
frame@f6eee000 = frame(4k)
frame@f6eef000 = frame(4k)
frame@f6ef0000 = frame(4k)
frame@f6ef1000 = frame(4k)
frame@f6ef2000 = frame(4k)
frame@f6ef3000 = frame(4k)
frame@f6ef4000 = frame(4k)
frame@f6ef5000 = frame(4k)
frame@f6ef6000 = frame(4k)
frame@f6ef7000 = frame(4k)
frame@f6ef8000 = frame(4k)
frame@f6ef9000 = frame(4k)
frame@f6efa000 = frame(4k)
frame@f6efb000 = frame(4k)
frame@f6efc000 = frame(4k)
frame@f6efd000 = frame(4k)
frame@f6efe000 = frame(4k)
frame@f6eff000 = frame(4k)
frame@f6f00000 = frame(4k)
frame@f6f01000 = frame(4k)
frame@f6f02000 = frame(4k)
frame@f6f03000 = frame(4k)
frame@f6f04000 = frame(4k)
frame@f6f05000 = frame(4k)
frame@f6f06000 = frame(4k)
frame@f6f07000 = frame(4k)
frame@f6f08000 = frame(4k)
frame@f6f09000 = frame(4k)
frame@f6f0a000 = frame(4k)
frame@f6f0b000 = frame(4k)
frame@f6f0c000 = frame(4k)
frame@f6f0d000 = frame(4k)
frame@f6f0e000 = frame(4k)
frame@f6f0f000 = frame(4k)
frame@f6f10000 = frame(4k)
frame@f6f11000 = frame(4k)
frame@f6f12000 = frame(4k)
frame@f6f13000 = frame(4k)
frame@f6f14000 = frame(4k)
frame@f6f15000 = frame(4k)
frame@f6f16000 = frame(4k)
frame@f6f17000 = frame(4k)
frame@f6f18000 = frame(4k)
frame@f6f19000 = frame(4k)
frame@f6f1a000 = frame(4k)
frame@f6f1b000 = frame(4k)
frame@f6f1c000 = frame(4k)
frame@f6f1d000 = frame(4k)
frame@f6f1e000 = frame(4k)
frame@f6f1f000 = frame(4k)
frame@f6f20000 = frame(4k)
frame@f6f21000 = frame(4k)
frame@f6f22000 = frame(4k)
frame@f6f23000 = frame(4k)
frame@f6f24000 = frame(4k)
frame@f6f25000 = frame(4k)
frame@f6f26000 = frame(4k)
frame@f6f27000 = frame(4k)
frame@f6f28000 = frame(4k)
frame@f6f29000 = frame(4k)
frame@f6f2a000 = frame(4k)
frame@f6f2b000 = frame(4k)
frame@f6f2c000 = frame(4k)
frame@f6f2d000 = frame(4k)
frame@f6f2e000 = frame(4k)
frame@f6f2f000 = frame(4k)
frame@f6f30000 = frame(4k)
frame@f6f31000 = frame(4k)
frame@f6f32000 = frame(4k)
frame@f6f33000 = frame(4k)
frame@f6f34000 = frame(4k)
frame@f6f35000 = frame(4k)
frame@f6f36000 = frame(4k)
frame@f6f37000 = frame(4k)
frame@f6f38000 = frame(4k)
frame@f6f39000 = frame(4k)
frame@f6f3a000 = frame(4k)
frame@f6f3b000 = frame(4k)
frame@f6f3c000 = frame(4k)
frame@f6f3d000 = frame(4k)
frame@f6f3e000 = frame(4k)
frame@f6f3f000 = frame(4k)
frame@f6f40000 = frame(4k)
frame@f6f41000 = frame(4k)
frame@f6f42000 = frame(4k)
frame@f6f43000 = frame(4k)
frame@f6f44000 = frame(4k)
frame@f6f45000 = frame(4k)
frame@f6f46000 = frame(4k)
frame@f6f47000 = frame(4k)
frame@f6f48000 = frame(4k)
frame@f6f49000 = frame(4k)
frame@f6f4a000 = frame(4k)
frame@f6f4b000 = frame(4k)
frame@f6f4c000 = frame(4k)
frame@f6f4d000 = frame(4k)
frame@f6f4e000 = frame(4k)
frame@f6f4f000 = frame(4k)
frame@f6f50000 = frame(4k)
frame@f6f51000 = frame(4k)
frame@f6f52000 = frame(4k)
frame@f6f53000 = frame(4k)
frame@f6f54000 = frame(4k)
frame@f6f55000 = frame(4k)
frame@f6f56000 = frame(4k)
frame@f6f57000 = frame(4k)
frame@f6f58000 = frame(4k)
frame@f6f59000 = frame(4k)
frame@f6f5a000 = frame(4k)
frame@f6f5b000 = frame(4k)
frame@f6f5c000 = frame(4k)
frame@f6f5d000 = frame(4k)
frame@f6f5e000 = frame(4k)
frame@f6f5f000 = frame(4k)
frame@f6f60000 = frame(4k)
frame@f6f61000 = frame(4k)
frame@f6f62000 = frame(4k)
frame@f6f63000 = frame(4k)
frame@f6f64000 = frame(4k)
frame@f6f65000 = frame(4k)
frame@f6f66000 = frame(4k)
frame@f6f67000 = frame(4k)
frame@f6f68000 = frame(4k)
frame@f6f69000 = frame(4k)
frame@f6f6a000 = frame(4k)
frame@f6f6b000 = frame(4k)
frame@f6f6c000 = frame(4k)
frame@f6f6d000 = frame(4k)
frame@f6f6e000 = frame(4k)
frame@f6f6f000 = frame(4k)
frame@f6f70000 = frame(4k)
frame@f6f71000 = frame(4k)
frame@f6f72000 = frame(4k)
frame@f6f73000 = frame(4k)
frame@f6f74000 = frame(4k)
frame@f6f75000 = frame(4k)
frame@f6f76000 = frame(4k)
frame@f6f77000 = frame(4k)
frame@f6f78000 = frame(4k)
frame@f6f79000 = frame(4k)
frame@f6f7a000 = frame(4k)
frame@f6f7b000 = frame(4k)
frame@f6f7c000 = frame(4k)
frame@f6f7d000 = frame(4k)
frame@f6f7e000 = frame(4k)
frame@f6f7f000 = frame(4k)
frame@f6f80000 = frame(4k)
frame@f6f81000 = frame(4k)
frame@f6f82000 = frame(4k)
frame@f6f83000 = frame(4k)
frame@f6f84000 = frame(4k)
frame@f6f85000 = frame(4k)
frame@f6f86000 = frame(4k)
frame@f6f87000 = frame(4k)
frame@f6f88000 = frame(4k)
frame@f6f89000 = frame(4k)
frame@f6f8a000 = frame(4k)
frame@f6f8b000 = frame(4k)
frame@f6f8c000 = frame(4k)
frame@f6f8d000 = frame(4k)
frame@f6f8e000 = frame(4k)
frame@f6f8f000 = frame(4k)
frame@f6f90000 = frame(4k)
frame@f6f91000 = frame(4k)
frame@f6f92000 = frame(4k)
frame@f6f93000 = frame(4k)
frame@f6f94000 = frame(4k)
frame@f6f95000 = frame(4k)
frame@f6f96000 = frame(4k)
frame@f6f97000 = frame(4k)
frame@f6f98000 = frame(4k)
frame@f6f99000 = frame(4k)
frame@f6f9a000 = frame(4k)
frame@f6f9b000 = frame(4k)
frame@f6f9c000 = frame(4k)
frame@f6f9d000 = frame(4k)
frame@f6f9e000 = frame(4k)
frame@f6f9f000 = frame(4k)
frame@f6fa0000 = frame(4k)
frame@f6fa1000 = frame(4k)
frame@f6fa2000 = frame(4k)
frame@f6fa3000 = frame(4k)
frame@f6fa4000 = frame(4k)
frame@f6fa5000 = frame(4k)
frame@f6fa6000 = frame(4k)
frame@f6fa7000 = frame(4k)
frame@f6fa8000 = frame(4k)
frame@f6fa9000 = frame(4k)
frame@f6faa000 = frame(4k)
frame@f6fab000 = frame(4k)
frame@f6fac000 = frame(4k)
frame@f6fad000 = frame(4k)
frame@f6fae000 = frame(4k)
frame@f6faf000 = frame(4k)
frame@f6fb0000 = frame(4k)
frame@f6fb1000 = frame(4k)
frame@f6fb2000 = frame(4k)
frame@f6fb3000 = frame(4k)
frame@f6fb4000 = frame(4k)
frame@f6fb5000 = frame(4k)
frame@f6fb6000 = frame(4k)
frame@f6fb7000 = frame(4k)
frame@f6fb8000 = frame(4k)
frame@f6fb9000 = frame(4k)
frame@f6fba000 = frame(4k)
frame@f6fbb000 = frame(4k)
frame@f6fbc000 = frame(4k)
frame@f6fbd000 = frame(4k)
frame@f6fbe000 = frame(4k)
frame@f6fbf000 = frame(4k)
frame@f6fc0000 = frame(4k)
frame@f6fc1000 = frame(4k)
frame@f6fc2000 = frame(4k)
frame@f6fc3000 = frame(4k)
frame@f6fc4000 = frame(4k)
frame@f6fc5000 = frame(4k)
frame@f6fc6000 = frame(4k)
frame@f6fc7000 = frame(4k)
frame@f6fc8000 = frame(4k)
frame@f6fc9000 = frame(4k)
frame@f6fca000 = frame(4k)
frame@f6fcb000 = frame(4k)
frame@f6fcc000 = frame(4k)
frame@f6fcd000 = frame(4k)
frame@f6fce000 = frame(4k)
frame@f6fcf000 = frame(4k)
frame@f6fd0000 = frame(4k)
frame@f6fd1000 = frame(4k)
frame@f6fd2000 = frame(4k)
frame@f6fd3000 = frame(4k)
frame@f6fd4000 = frame(4k)
frame@f6fd5000 = frame(4k)
frame@f6fd6000 = frame(4k)
frame@f6fd7000 = frame(4k)
frame@f6fd8000 = frame(4k)
frame@f6fd9000 = frame(4k)
frame@f6fda000 = frame(4k)
frame@f6fdb000 = frame(4k)
frame@f6fdc000 = frame(4k)
frame@f6fdd000 = frame(4k)
frame@f6fde000 = frame(4k)
frame@f6fdf000 = frame(4k)
frame@f6fe0000 = frame(4k)
frame@f6fe1000 = frame(4k)
frame@f6fe2000 = frame(4k)
frame@f6fe3000 = frame(4k)
frame@f6fe4000 = frame(4k)
frame@f6fe5000 = frame(4k)
frame@f6fe6000 = frame(4k)
frame@f6fe7000 = frame(4k)
frame@f6fe8000 = frame(4k)
frame@f6fe9000 = frame(4k)
frame@f6fea000 = frame(4k)
frame@f6feb000 = frame(4k)
frame@f6fec000 = frame(4k)
frame@f6fed000 = frame(4k)
frame@f6fee000 = frame(4k)
frame@f6fef000 = frame(4k)
frame@f6ff0000 = frame(4k)
frame@f6ff1000 = frame(4k)
frame@f6ff2000 = frame(4k)
frame@f6ff3000 = frame(4k)
frame@f6ff4000 = frame(4k)
frame@f6ff5000 = frame(4k)
frame@f6ff6000 = frame(4k)
frame@f6ff7000 = frame(4k)
frame@f6ff8000 = frame(4k)
frame@f6ff9000 = frame(4k)
frame@f6ffa000 = frame(4k)
frame@f6ffb000 = frame(4k)
frame@f6ffc000 = frame(4k)
frame@f6ffd000 = frame(4k)
frame@f6ffe000 = frame(4k)
frame@f6fff000 = frame(4k)
frame@f7000000 = frame(4k)
frame@f7001000 = frame(4k)
frame@f7002000 = frame(4k)
frame@f7003000 = frame(4k)
frame@f7004000 = frame(4k)
frame@f7005000 = frame(4k)
frame@f7006000 = frame(4k)
frame@f7007000 = frame(4k)
frame@f7008000 = frame(4k)
frame@f7009000 = frame(4k)
frame@f700a000 = frame(4k)
frame@f700b000 = frame(4k)
frame@f700c000 = frame(4k)
frame@f700d000 = frame(4k)
frame@f700e000 = frame(4k)
frame@f700f000 = frame(4k)
frame@f7010000 = frame(4k)
frame@f7011000 = frame(4k)
frame@f7012000 = frame(4k)
frame@f7013000 = frame(4k)
frame@f7014000 = frame(4k)
frame@f7015000 = frame(4k)
frame@f7016000 = frame(4k)
frame@f7017000 = frame(4k)
frame@f7018000 = frame(4k)
frame@f7019000 = frame(4k)
frame@f701a000 = frame(4k)
frame@f701b000 = frame(4k)
frame@f701c000 = frame(4k)
frame@f701d000 = frame(4k)
frame@f701e000 = frame(4k)
frame@f701f000 = frame(4k)
frame@f7020000 = frame(4k)
frame@f7021000 = frame(4k)
frame@f7022000 = frame(4k)
frame@f7023000 = frame(4k)
frame@f7024000 = frame(4k)
frame@f7025000 = frame(4k)
frame@f7026000 = frame(4k)
frame@f7027000 = frame(4k)
frame@f7028000 = frame(4k)
frame@f7029000 = frame(4k)
frame@f702a000 = frame(4k)
frame@f702b000 = frame(4k)
frame@f702c000 = frame(4k)
frame@f702d000 = frame(4k)
frame@f702e000 = frame(4k)
frame@f702f000 = frame(4k)
frame@f7030000 = frame(4k)
frame@f7031000 = frame(4k)
frame@f7032000 = frame(4k)
frame@f7033000 = frame(4k)
frame@f7034000 = frame(4k)
frame@f7035000 = frame(4k)
frame@f7036000 = frame(4k)
frame@f7037000 = frame(4k)
frame@f7038000 = frame(4k)
frame@f7039000 = frame(4k)
frame@f703a000 = frame(4k)
frame@f703b000 = frame(4k)
frame@f703c000 = frame(4k)
frame@f703d000 = frame(4k)
frame@f703e000 = frame(4k)
frame@f703f000 = frame(4k)
frame@f7040000 = frame(4k)
frame@f7041000 = frame(4k)
frame@f7042000 = frame(4k)
frame@f7043000 = frame(4k)
frame@f7044000 = frame(4k)
frame@f7045000 = frame(4k)
frame@f7046000 = frame(4k)
frame@f7047000 = frame(4k)
frame@f7048000 = frame(4k)
frame@f7049000 = frame(4k)
frame@f704a000 = frame(4k)
frame@f704b000 = frame(4k)
frame@f704c000 = frame(4k)
frame@f704d000 = frame(4k)
frame@f704e000 = frame(4k)
frame@f704f000 = frame(4k)
frame@f7050000 = frame(4k)
frame@f7051000 = frame(4k)
frame@f7052000 = frame(4k)
frame@f7053000 = frame(4k)
frame@f7054000 = frame(4k)
frame@f7055000 = frame(4k)
frame@f7056000 = frame(4k)
frame@f7057000 = frame(4k)
frame@f7058000 = frame(4k)
frame@f7059000 = frame(4k)
frame@f705a000 = frame(4k)
frame@f705b000 = frame(4k)
frame@f705c000 = frame(4k)
frame@f705d000 = frame(4k)
frame@f705e000 = frame(4k)
frame@f705f000 = frame(4k)
frame@f7060000 = frame(4k)
frame@f7061000 = frame(4k)
frame@f7062000 = frame(4k)
frame@f7063000 = frame(4k)
frame@f7064000 = frame(4k)
frame@f7065000 = frame(4k)
frame@f7066000 = frame(4k)
frame@f7067000 = frame(4k)
frame@f7068000 = frame(4k)
frame@f7069000 = frame(4k)
frame@f706a000 = frame(4k)
frame@f706b000 = frame(4k)
frame@f706c000 = frame(4k)
frame@f706d000 = frame(4k)
frame@f706e000 = frame(4k)
frame@f706f000 = frame(4k)
frame@f7070000 = frame(4k)
frame@f7071000 = frame(4k)
frame@f7072000 = frame(4k)
frame@f7073000 = frame(4k)
frame@f7074000 = frame(4k)
frame@f7075000 = frame(4k)
frame@f7076000 = frame(4k)
frame@f7077000 = frame(4k)
frame@f7078000 = frame(4k)
frame@f7079000 = frame(4k)
frame@f707a000 = frame(4k)
frame@f707b000 = frame(4k)
frame@f707c000 = frame(4k)
frame@f707d000 = frame(4k)
frame@f707e000 = frame(4k)
frame@f707f000 = frame(4k)
frame@f7080000 = frame(4k)
frame@f7081000 = frame(4k)
frame@f7082000 = frame(4k)
frame@f7083000 = frame(4k)
frame@f7084000 = frame(4k)
frame@f7085000 = frame(4k)
frame@f7086000 = frame(4k)
frame@f7087000 = frame(4k)
frame@f7088000 = frame(4k)
frame@f7089000 = frame(4k)
frame@f708a000 = frame(4k)
frame@f708b000 = frame(4k)
frame@f708c000 = frame(4k)
frame@f708d000 = frame(4k)
frame@f708e000 = frame(4k)
frame@f708f000 = frame(4k)
frame@f7090000 = frame(4k)
frame@f7091000 = frame(4k)
frame@f7092000 = frame(4k)
frame@f7093000 = frame(4k)
frame@f7094000 = frame(4k)
frame@f7095000 = frame(4k)
frame@f7096000 = frame(4k)
frame@f7097000 = frame(4k)
frame@f7098000 = frame(4k)
frame@f7099000 = frame(4k)
frame@f709a000 = frame(4k)
frame@f709b000 = frame(4k)
frame@f709c000 = frame(4k)
frame@f709d000 = frame(4k)
frame@f709e000 = frame(4k)
frame@f709f000 = frame(4k)
frame@f70a0000 = frame(4k)
frame@f70a1000 = frame(4k)
frame@f70a2000 = frame(4k)
frame@f70a3000 = frame(4k)
frame@f70a4000 = frame(4k)
frame@f70a5000 = frame(4k)
frame@f70a6000 = frame(4k)
frame@f70a7000 = frame(4k)
frame@f70a8000 = frame(4k)
frame@f70a9000 = frame(4k)
frame@f70aa000 = frame(4k)
frame@f70ab000 = frame(4k)
frame@f70ac000 = frame(4k)
frame@f70ad000 = frame(4k)
frame@f70ae000 = frame(4k)
frame@f70af000 = frame(4k)
frame@f70b0000 = frame(4k)
frame@f70b1000 = frame(4k)
frame@f70b2000 = frame(4k)
frame@f70b3000 = frame(4k)
frame@f70b4000 = frame(4k)
frame@f70b5000 = frame(4k)
frame@f70b6000 = frame(4k)
frame@f70b7000 = frame(4k)
frame@f70b8000 = frame(4k)
frame@f70b9000 = frame(4k)
frame@f70ba000 = frame(4k)
frame@f70bb000 = frame(4k)
frame@f70bc000 = frame(4k)
frame@f70bd000 = frame(4k)
frame@f70be000 = frame(4k)
frame@f70bf000 = frame(4k)
frame@f70c0000 = frame(4k)
frame@f70c1000 = frame(4k)
frame@f70c2000 = frame(4k)
frame@f70c3000 = frame(4k)
frame@f70c4000 = frame(4k)
frame@f70c5000 = frame(4k)
frame@f70c6000 = frame(4k)
frame@f70c7000 = frame(4k)
frame@f70c8000 = frame(4k)
frame@f70c9000 = frame(4k)
frame@f70ca000 = frame(4k)
frame@f70cb000 = frame(4k)
frame@f70cc000 = frame(4k)
frame@f70cd000 = frame(4k)
frame@f70ce000 = frame(4k)
frame@f70cf000 = frame(4k)
frame@f70d0000 = frame(4k)
frame@f70d1000 = frame(4k)
frame@f70d2000 = frame(4k)
frame@f70d3000 = frame(4k)
frame@f70d4000 = frame(4k)
frame@f70d5000 = frame(4k)
frame@f70d6000 = frame(4k)
frame@f70d7000 = frame(4k)
frame@f70d8000 = frame(4k)
frame@f70d9000 = frame(4k)
frame@f70da000 = frame(4k)
frame@f70db000 = frame(4k)
frame@f70dc000 = frame(4k)
frame@f70dd000 = frame(4k)
frame@f70de000 = frame(4k)
frame@f70df000 = frame(4k)
frame@f70e0000 = frame(4k)
frame@f70e1000 = frame(4k)
frame@f70e2000 = frame(4k)
frame@f70e3000 = frame(4k)
frame@f70e4000 = frame(4k)
frame@f70e5000 = frame(4k)
frame@f70e6000 = frame(4k)
frame@f70e7000 = frame(4k)
frame@f70e8000 = frame(4k)
frame@f70e9000 = frame(4k)
frame@f70ea000 = frame(4k)
frame@f70eb000 = frame(4k)
frame@f70ec000 = frame(4k)
frame@f70ed000 = frame(4k)
frame@f70ee000 = frame(4k)
frame@f70ef000 = frame(4k)
frame@f70f0000 = frame(4k)
frame@f70f1000 = frame(4k)
frame@f70f2000 = frame(4k)
frame@f70f3000 = frame(4k)
frame@f70f4000 = frame(4k)
frame@f70f5000 = frame(4k)
frame@f70f6000 = frame(4k)
frame@f70f7000 = frame(4k)
frame@f70f8000 = frame(4k)
frame@f70f9000 = frame(4k)
frame@f70fa000 = frame(4k)
frame@f70fb000 = frame(4k)
frame@f70fc000 = frame(4k)
frame@f70fd000 = frame(4k)
frame@f70fe000 = frame(4k)
frame@f70ff000 = frame(4k)
frame@f7100000 = frame(4k)
frame@f7101000 = frame(4k)
frame@f7102000 = frame(4k)
frame@f7103000 = frame(4k)
frame@f7104000 = frame(4k)
frame@f7105000 = frame(4k)
frame@f7106000 = frame(4k)
frame@f7107000 = frame(4k)
frame@f7108000 = frame(4k)
frame@f7109000 = frame(4k)
frame@f710a000 = frame(4k)
frame@f710b000 = frame(4k)
frame@f710c000 = frame(4k)
frame@f710d000 = frame(4k)
frame@f710e000 = frame(4k)
frame@f710f000 = frame(4k)
frame@f7110000 = frame(4k)
frame@f7111000 = frame(4k)
frame@f7112000 = frame(4k)
frame@f7113000 = frame(4k)
frame@f7114000 = frame(4k)
frame@f7115000 = frame(4k)
frame@f7116000 = frame(4k)
frame@f7117000 = frame(4k)
frame@f7118000 = frame(4k)
frame@f7119000 = frame(4k)
frame@f711a000 = frame(4k)
frame@f711b000 = frame(4k)
frame@f711c000 = frame(4k)
frame@f711d000 = frame(4k)
frame@f711e000 = frame(4k)
frame@f711f000 = frame(4k)
frame@f7120000 = frame(4k)
frame@f7121000 = frame(4k)
frame@f7122000 = frame(4k)
frame@f7123000 = frame(4k)
frame@f7124000 = frame(4k)
frame@f7125000 = frame(4k)
frame@f7126000 = frame(4k)
frame@f7127000 = frame(4k)
frame@f7128000 = frame(4k)
frame@f7129000 = frame(4k)
frame@f712a000 = frame(4k)
frame@f712b000 = frame(4k)
frame@f712c000 = frame(4k)
frame@f712d000 = frame(4k)
frame@f712e000 = frame(4k)
frame@f712f000 = frame(4k)
frame@f7130000 = frame(4k)
frame@f7131000 = frame(4k)
frame@f7132000 = frame(4k)
frame@f7133000 = frame(4k)
frame@f7134000 = frame(4k)
frame@f7135000 = frame(4k)
frame@f7136000 = frame(4k)
frame@f7137000 = frame(4k)
frame@f7138000 = frame(4k)
frame@f7139000 = frame(4k)
frame@f713a000 = frame(4k)
frame@f713b000 = frame(4k)
frame@f713c000 = frame(4k)
frame@f713d000 = frame(4k)
frame@f713e000 = frame(4k)
frame@f713f000 = frame(4k)
frame@f7140000 = frame(4k)
frame@f7141000 = frame(4k)
frame@f7142000 = frame(4k)
frame@f7143000 = frame(4k)
frame@f7144000 = frame(4k)
frame@f7145000 = frame(4k)
frame@f7146000 = frame(4k)
frame@f7147000 = frame(4k)
frame@f7148000 = frame(4k)
frame@f7149000 = frame(4k)
frame@f714a000 = frame(4k)
frame@f714b000 = frame(4k)
frame@f714c000 = frame(4k)
frame@f714d000 = frame(4k)
frame@f714e000 = frame(4k)
frame@f714f000 = frame(4k)
frame@f7150000 = frame(4k)
frame@f7151000 = frame(4k)
frame@f7152000 = frame(4k)
frame@f7153000 = frame(4k)
frame@f7154000 = frame(4k)
frame@f7155000 = frame(4k)
frame@f7156000 = frame(4k)
frame@f7157000 = frame(4k)
frame@f7158000 = frame(4k)
frame@f7159000 = frame(4k)
frame@f715a000 = frame(4k)
frame@f715b000 = frame(4k)
frame@f715c000 = frame(4k)
frame@f715d000 = frame(4k)
frame@f715e000 = frame(4k)
frame@f715f000 = frame(4k)
frame@f7160000 = frame(4k)
frame@f7161000 = frame(4k)
frame@f7162000 = frame(4k)
frame@f7163000 = frame(4k)
frame@f7164000 = frame(4k)
frame@f7165000 = frame(4k)
frame@f7166000 = frame(4k)
frame@f7167000 = frame(4k)
frame@f7168000 = frame(4k)
frame@f7169000 = frame(4k)
frame@f716a000 = frame(4k)
frame@f716b000 = frame(4k)
frame@f716c000 = frame(4k)
frame@f716d000 = frame(4k)
frame@f716e000 = frame(4k)
frame@f716f000 = frame(4k)
frame@f7170000 = frame(4k)
frame@f7171000 = frame(4k)
frame@f7172000 = frame(4k)
frame@f7173000 = frame(4k)
frame@f7174000 = frame(4k)
frame@f7175000 = frame(4k)
frame@f7176000 = frame(4k)
frame@f7177000 = frame(4k)
frame@f7178000 = frame(4k)
frame@f7179000 = frame(4k)
frame@f717a000 = frame(4k)
frame@f717b000 = frame(4k)
frame@f717c000 = frame(4k)
frame@f717d000 = frame(4k)
frame@f717e000 = frame(4k)
frame@f717f000 = frame(4k)
frame@f7180000 = frame(4k)
frame@f7181000 = frame(4k)
frame@f7182000 = frame(4k)
frame@f7183000 = frame(4k)
frame@f7184000 = frame(4k)
frame@f7185000 = frame(4k)
frame@f7186000 = frame(4k)
frame@f7187000 = frame(4k)
frame@f7188000 = frame(4k)
frame@f7189000 = frame(4k)
frame@f718a000 = frame(4k)
frame@f718b000 = frame(4k)
frame@f718c000 = frame(4k)
frame@f718d000 = frame(4k)
frame@f718e000 = frame(4k)
frame@f718f000 = frame(4k)
frame@f7190000 = frame(4k)
frame@f7191000 = frame(4k)
frame@f7192000 = frame(4k)
frame@f7193000 = frame(4k)
frame@f7194000 = frame(4k)
frame@f7195000 = frame(4k)
frame@f7196000 = frame(4k)
frame@f7197000 = frame(4k)
frame@f7198000 = frame(4k)
frame@f7199000 = frame(4k)
frame@f719a000 = frame(4k)
frame@f719b000 = frame(4k)
frame@f719c000 = frame(4k)
frame@f719d000 = frame(4k)
frame@f719e000 = frame(4k)
frame@f719f000 = frame(4k)
frame@f71a0000 = frame(4k)
frame@f71a1000 = frame(4k)
frame@f71a2000 = frame(4k)
frame@f71a3000 = frame(4k)
frame@f71a4000 = frame(4k)
frame@f71a5000 = frame(4k)
frame@f71a6000 = frame(4k)
frame@f71a7000 = frame(4k)
frame@f71a8000 = frame(4k)
frame@f71a9000 = frame(4k)
frame@f71aa000 = frame(4k)
frame@f71ab000 = frame(4k)
frame@f71ac000 = frame(4k)
frame@f71ad000 = frame(4k)
frame@f71ae000 = frame(4k)
frame@f71af000 = frame(4k)
frame@f71b0000 = frame(4k)
frame@f71b1000 = frame(4k)
frame@f71b2000 = frame(4k)
frame@f71b3000 = frame(4k)
frame@f71b4000 = frame(4k)
frame@f71b5000 = frame(4k)
frame@f71b6000 = frame(4k)
frame@f71b7000 = frame(4k)
frame@f71b8000 = frame(4k)
frame@f71b9000 = frame(4k)
frame@f71ba000 = frame(4k)
frame@f71bb000 = frame(4k)
frame@f71bc000 = frame(4k)
frame@f71bd000 = frame(4k)
frame@f71be000 = frame(4k)
frame@f71bf000 = frame(4k)
frame@f71c0000 = frame(4k)
frame@f71c1000 = frame(4k)
frame@f71c2000 = frame(4k)
frame@f71c3000 = frame(4k)
frame@f71c4000 = frame(4k)
frame@f71c5000 = frame(4k)
frame@f71c6000 = frame(4k)
frame@f71c7000 = frame(4k)
frame@f71c8000 = frame(4k)
frame@f71c9000 = frame(4k)
frame@f71ca000 = frame(4k)
frame@f71cb000 = frame(4k)
frame@f71cc000 = frame(4k)
frame@f71cd000 = frame(4k)
frame@f71ce000 = frame(4k)
frame@f71cf000 = frame(4k)
frame@f71d0000 = frame(4k)
frame@f71d1000 = frame(4k)
frame@f71d2000 = frame(4k)
frame@f71d3000 = frame(4k)
frame@f71d4000 = frame(4k)
frame@f71d5000 = frame(4k)
frame@f71d6000 = frame(4k)
frame@f71d7000 = frame(4k)
frame@f71d8000 = frame(4k)
frame@f71d9000 = frame(4k)
frame@f71da000 = frame(4k)
frame@f71db000 = frame(4k)
frame@f71dc000 = frame(4k)
frame@f71dd000 = frame(4k)
frame@f71de000 = frame(4k)
frame@f71df000 = frame(4k)
frame@f71e0000 = frame(4k)
frame@f71e1000 = frame(4k)
frame@f71e2000 = frame(4k)
frame@f71e3000 = frame(4k)
frame@f71e4000 = frame(4k)
frame@f71e5000 = frame(4k)
frame@f71e6000 = frame(4k)
frame@f71e7000 = frame(4k)
frame@f71e8000 = frame(4k)
frame@f71e9000 = frame(4k)
frame@f71ea000 = frame(4k)
frame@f71eb000 = frame(4k)
frame@f71ec000 = frame(4k)
frame@f71ed000 = frame(4k)
frame@f71ee000 = frame(4k)
frame@f71ef000 = frame(4k)
frame@f71f0000 = frame(4k)
frame@f71f1000 = frame(4k)
frame@f71f2000 = frame(4k)
frame@f71f3000 = frame(4k)
frame@f71f4000 = frame(4k)
frame@f71f5000 = frame(4k)
frame@f71f6000 = frame(4k)
frame@f71f7000 = frame(4k)
frame@f71f8000 = frame(4k)
frame@f71f9000 = frame(4k)
frame@f71fa000 = frame(4k)
frame@f71fb000 = frame(4k)
frame@f71fc000 = frame(4k)
frame@f71fd000 = frame(4k)
frame@f71fe000 = frame(4k)
frame@f71ff000 = frame(4k)
frame@f7200000 = frame(4k)
frame@f7201000 = frame(4k)
frame@f7202000 = frame(4k)
frame@f7203000 = frame(4k)
frame@f7204000 = frame(4k)
frame@f7205000 = frame(4k)
frame@f7206000 = frame(4k)
frame@f7207000 = frame(4k)
frame@f7208000 = frame(4k)
frame@f7209000 = frame(4k)
frame@f720a000 = frame(4k)
frame@f720b000 = frame(4k)
frame@f720c000 = frame(4k)
frame@f720d000 = frame(4k)
frame@f720e000 = frame(4k)
frame@f720f000 = frame(4k)
frame@f7210000 = frame(4k)
frame@f7211000 = frame(4k)
frame@f7212000 = frame(4k)
frame@f7213000 = frame(4k)
frame@f7214000 = frame(4k)
frame@f7215000 = frame(4k)
frame@f7216000 = frame(4k)
frame@f7217000 = frame(4k)
frame@f7218000 = frame(4k)
frame@f7219000 = frame(4k)
frame@f721a000 = frame(4k)
frame@f721b000 = frame(4k)
frame@f721c000 = frame(4k)
frame@f721d000 = frame(4k)
frame@f721e000 = frame(4k)
frame@f721f000 = frame(4k)
frame@f7220000 = frame(4k)
frame@f7221000 = frame(4k)
frame@f7222000 = frame(4k)
frame@f7223000 = frame(4k)
frame@f7224000 = frame(4k)
frame@f7225000 = frame(4k)
frame@f7226000 = frame(4k)
frame@f7227000 = frame(4k)
frame@f7228000 = frame(4k)
frame@f7229000 = frame(4k)
frame@f722a000 = frame(4k)
frame@f722b000 = frame(4k)
frame@f722c000 = frame(4k)
frame@f722d000 = frame(4k)
frame@f722e000 = frame(4k)
frame@f722f000 = frame(4k)
frame@f7230000 = frame(4k)
frame@f7231000 = frame(4k)
frame@f7232000 = frame(4k)
frame@f7233000 = frame(4k)
frame@f7234000 = frame(4k)
frame@f7235000 = frame(4k)
frame@f7236000 = frame(4k)
frame@f7237000 = frame(4k)
frame@f7238000 = frame(4k)
frame@f7239000 = frame(4k)
frame@f723a000 = frame(4k)
frame@f723b000 = frame(4k)
frame@f723c000 = frame(4k)
frame@f723d000 = frame(4k)
frame@f723e000 = frame(4k)
frame@f723f000 = frame(4k)
frame@f7240000 = frame(4k)
frame@f7241000 = frame(4k)
frame@f7242000 = frame(4k)
frame@f7243000 = frame(4k)
frame@f7244000 = frame(4k)
frame@f7245000 = frame(4k)
frame@f7246000 = frame(4k)
frame@f7247000 = frame(4k)
frame@f7248000 = frame(4k)
frame@f7249000 = frame(4k)
frame@f724a000 = frame(4k)
frame@f724b000 = frame(4k)
frame@f724c000 = frame(4k)
frame@f724d000 = frame(4k)
frame@f724e000 = frame(4k)
frame@f724f000 = frame(4k)
frame@f7250000 = frame(4k)
frame@f7251000 = frame(4k)
frame@f7252000 = frame(4k)
frame@f7253000 = frame(4k)
frame@f7254000 = frame(4k)
frame@f7255000 = frame(4k)
frame@f7256000 = frame(4k)
frame@f7257000 = frame(4k)
frame@f7258000 = frame(4k)
frame@f7259000 = frame(4k)
frame@f725a000 = frame(4k)
frame@f725b000 = frame(4k)
frame@f725c000 = frame(4k)
frame@f725d000 = frame(4k)
frame@f725e000 = frame(4k)
frame@f725f000 = frame(4k)
frame@f7260000 = frame(4k)
frame@f7261000 = frame(4k)
frame@f7262000 = frame(4k)
frame@f7263000 = frame(4k)
frame@f7264000 = frame(4k)
frame@f7265000 = frame(4k)
frame@f7266000 = frame(4k)
frame@f7267000 = frame(4k)
frame@f7268000 = frame(4k)
frame@f7269000 = frame(4k)
frame@f726a000 = frame(4k)
frame@f726b000 = frame(4k)
frame@f726c000 = frame(4k)
frame@f726d000 = frame(4k)
frame@f726e000 = frame(4k)
frame@f726f000 = frame(4k)
frame@f7270000 = frame(4k)
frame@f7271000 = frame(4k)
frame@f7272000 = frame(4k)
frame@f7273000 = frame(4k)
frame@f7274000 = frame(4k)
frame@f7275000 = frame(4k)
frame@f7276000 = frame(4k)
frame@f7277000 = frame(4k)
frame@f7278000 = frame(4k)
frame@f7279000 = frame(4k)
frame@f727a000 = frame(4k)
frame@f727b000 = frame(4k)
frame@f727c000 = frame(4k)
frame@f727d000 = frame(4k)
frame@f727e000 = frame(4k)
frame@f727f000 = frame(4k)
frame@f7280000 = frame(4k)
frame@f7281000 = frame(4k)
frame@f7282000 = frame(4k)
frame@f7283000 = frame(4k)
frame@f7284000 = frame(4k)
frame@f7285000 = frame(4k)
frame@f7286000 = frame(4k)
frame@f7287000 = frame(4k)
frame@f7288000 = frame(4k)
frame@f7289000 = frame(4k)
frame@f728a000 = frame(4k)
frame@f728b000 = frame(4k)
frame@f728c000 = frame(4k)
frame@f728d000 = frame(4k)
frame@f728e000 = frame(4k)
frame@f728f000 = frame(4k)
frame@f7290000 = frame(4k)
frame@f7291000 = frame(4k)
frame@f7292000 = frame(4k)
frame@f7293000 = frame(4k)
frame@f7294000 = frame(4k)
frame@f7295000 = frame(4k)
frame@f7296000 = frame(4k)
frame@f7297000 = frame(4k)
frame@f7298000 = frame(4k)
frame@f7299000 = frame(4k)
frame@f729a000 = frame(4k)
frame@f729b000 = frame(4k)
frame@f729c000 = frame(4k)
frame@f729d000 = frame(4k)
frame@f729e000 = frame(4k)
frame@f729f000 = frame(4k)
frame@f72a0000 = frame(4k)
frame@f72a1000 = frame(4k)
frame@f72a2000 = frame(4k)
frame@f72a3000 = frame(4k)
frame@f72a4000 = frame(4k)
frame@f72a5000 = frame(4k)
frame@f72a6000 = frame(4k)
frame@f72a7000 = frame(4k)
frame@f72a8000 = frame(4k)
frame@f72a9000 = frame(4k)
frame@f72aa000 = frame(4k)
frame@f72ab000 = frame(4k)
frame@f72ac000 = frame(4k)
frame@f72ad000 = frame(4k)
frame@f72ae000 = frame(4k)
frame@f72af000 = frame(4k)
frame@f72b0000 = frame(4k)
frame@f72b1000 = frame(4k)
frame@f72b2000 = frame(4k)
frame@f72b3000 = frame(4k)
frame@f72b4000 = frame(4k)
frame@f72b5000 = frame(4k)
frame@f72b6000 = frame(4k)
frame@f72b7000 = frame(4k)
frame@f72b8000 = frame(4k)
frame@f72b9000 = frame(4k)
frame@f72ba000 = frame(4k)
frame@f72bb000 = frame(4k)
frame@f72bc000 = frame(4k)
frame@f72bd000 = frame(4k)
frame@f72be000 = frame(4k)
frame@f72bf000 = frame(4k)
frame@f72c0000 = frame(4k)
frame@f72c1000 = frame(4k)
frame@f72c2000 = frame(4k)
frame@f72c3000 = frame(4k)
frame@f72c4000 = frame(4k)
frame@f72c5000 = frame(4k)
frame@f72c6000 = frame(4k)
frame@f72c7000 = frame(4k)
frame@f72c8000 = frame(4k)
frame@f72c9000 = frame(4k)
frame@f72ca000 = frame(4k)
frame@f72cb000 = frame(4k)
frame@f72cc000 = frame(4k)
frame@f72cd000 = frame(4k)
frame@f72ce000 = frame(4k)
frame@f72cf000 = frame(4k)
frame@f72d0000 = frame(4k)
frame@f72d1000 = frame(4k)
frame@f72d2000 = frame(4k)
frame@f72d3000 = frame(4k)
frame@f72d4000 = frame(4k)
frame@f72d5000 = frame(4k)
frame@f72d6000 = frame(4k)
frame@f72d7000 = frame(4k)
frame@f72d8000 = frame(4k)
frame@f72d9000 = frame(4k)
frame@f72da000 = frame(4k)
frame@f72db000 = frame(4k)
frame@f72dc000 = frame(4k)
frame@f72dd000 = frame(4k)
frame@f72de000 = frame(4k)
frame@f72df000 = frame(4k)
frame@f72e0000 = frame(4k)
frame@f72e1000 = frame(4k)
frame@f72e2000 = frame(4k)
frame@f72e3000 = frame(4k)
frame@f72e4000 = frame(4k)
frame@f72e5000 = frame(4k)
frame@f72e6000 = frame(4k)
frame@f72e7000 = frame(4k)
frame@f72e8000 = frame(4k)
frame@f72e9000 = frame(4k)
frame@f72ea000 = frame(4k)
frame@f72eb000 = frame(4k)
frame@f72ec000 = frame(4k)
frame@f72ed000 = frame(4k)
frame@f72ee000 = frame(4k)
frame@f72ef000 = frame(4k)
frame@f72f0000 = frame(4k)
frame@f72f1000 = frame(4k)
frame@f72f2000 = frame(4k)
frame@f72f3000 = frame(4k)
frame@f72f4000 = frame(4k)
frame@f72f5000 = frame(4k)
frame@f72f6000 = frame(4k)
frame@f72f7000 = frame(4k)
frame@f72f8000 = frame(4k)
frame@f72f9000 = frame(4k)
frame@f72fa000 = frame(4k)
frame@f72fb000 = frame(4k)
frame@f72fc000 = frame(4k)
frame@f72fd000 = frame(4k)
frame@f72fe000 = frame(4k)
frame@f72ff000 = frame(4k)
frame@f9800000 = frame(4k)
frame@f9801000 = frame(4k)
frame@f9802000 = frame(4k)
frame@f9803000 = frame(4k)
frame@f9804000 = frame(4k)
frame@f9805000 = frame(4k)
frame@f9806000 = frame(4k)
frame@f9807000 = frame(4k)
frame@f9808000 = frame(4k)
frame@f9809000 = frame(4k)
frame@f980a000 = frame(4k)
frame@f980b000 = frame(4k)
frame@f980c000 = frame(4k)
frame@f980d000 = frame(4k)
frame@f980e000 = frame(4k)
frame@f980f000 = frame(4k)
frame@f9810000 = frame(4k)
frame@f9811000 = frame(4k)
frame@f9812000 = frame(4k)
frame@f9813000 = frame(4k)
frame@f9814000 = frame(4k)
frame@f9815000 = frame(4k)
frame@f9816000 = frame(4k)
frame@f9817000 = frame(4k)
frame@f9818000 = frame(4k)
frame@f9819000 = frame(4k)
frame@f981a000 = frame(4k)
frame@f981b000 = frame(4k)
frame@f981c000 = frame(4k)
frame@f981d000 = frame(4k)
frame@f981e000 = frame(4k)
frame@f981f000 = frame(4k)
frame@f9820000 = frame(4k)
frame@f9821000 = frame(4k)
frame@f9822000 = frame(4k)
frame@f9823000 = frame(4k)
frame@f9824000 = frame(4k)
frame@f9825000 = frame(4k)
frame@f9826000 = frame(4k)
frame@f9827000 = frame(4k)
frame@f9828000 = frame(4k)
frame@f9829000 = frame(4k)
frame@f982a000 = frame(4k)
frame@f982b000 = frame(4k)
frame@f982c000 = frame(4k)
frame@f982d000 = frame(4k)
frame@f982e000 = frame(4k)
frame@f982f000 = frame(4k)
frame@f9830000 = frame(4k)
frame@f9831000 = frame(4k)
frame@f9832000 = frame(4k)
frame@f9833000 = frame(4k)
frame@f9834000 = frame(4k)
frame@f9835000 = frame(4k)
frame@f9836000 = frame(4k)
frame@f9837000 = frame(4k)
frame@f9838000 = frame(4k)
frame@f9839000 = frame(4k)
frame@f983a000 = frame(4k)
frame@f983b000 = frame(4k)
frame@f983c000 = frame(4k)
frame@f983d000 = frame(4k)
frame@f983e000 = frame(4k)
frame@f983f000 = frame(4k)
frame@f9840000 = frame(4k)
frame@f9841000 = frame(4k)
frame@f9842000 = frame(4k)
frame@f9843000 = frame(4k)
frame@f9844000 = frame(4k)
frame@f9845000 = frame(4k)
frame@f9846000 = frame(4k)
frame@f9847000 = frame(4k)
frame@f9848000 = frame(4k)
frame@f9849000 = frame(4k)
frame@f984a000 = frame(4k)
frame@f984b000 = frame(4k)
frame@f984c000 = frame(4k)
frame@f984d000 = frame(4k)
frame@f984e000 = frame(4k)
frame@f984f000 = frame(4k)
frame@f9850000 = frame(4k)
frame@f9851000 = frame(4k)
frame@f9852000 = frame(4k)
frame@f9853000 = frame(4k)
frame@f9854000 = frame(4k)
frame@f9855000 = frame(4k)
frame@f9856000 = frame(4k)
frame@f9857000 = frame(4k)
frame@f9858000 = frame(4k)
frame@f9859000 = frame(4k)
frame@f985a000 = frame(4k)
frame@f985b000 = frame(4k)
frame@f985c000 = frame(4k)
frame@f985d000 = frame(4k)
frame@f985e000 = frame(4k)
frame@f985f000 = frame(4k)
frame@f9860000 = frame(4k)
frame@f9861000 = frame(4k)
frame@f9862000 = frame(4k)
frame@f9863000 = frame(4k)
frame@f9864000 = frame(4k)
frame@f9865000 = frame(4k)
frame@f9866000 = frame(4k)
frame@f9867000 = frame(4k)
frame@f9868000 = frame(4k)
frame@f9869000 = frame(4k)
frame@f986a000 = frame(4k)
frame@f986b000 = frame(4k)
frame@f986c000 = frame(4k)
frame@f986d000 = frame(4k)
frame@f986e000 = frame(4k)
frame@f986f000 = frame(4k)
frame@f9870000 = frame(4k)
frame@f9871000 = frame(4k)
frame@f9872000 = frame(4k)
frame@f9873000 = frame(4k)
frame@f9874000 = frame(4k)
frame@f9875000 = frame(4k)
frame@f9876000 = frame(4k)
frame@f9877000 = frame(4k)
frame@f9878000 = frame(4k)
frame@f9879000 = frame(4k)
frame@f987a000 = frame(4k)
frame@f987b000 = frame(4k)
frame@f987c000 = frame(4k)
frame@f987d000 = frame(4k)
frame@f987e000 = frame(4k)
frame@f987f000 = frame(4k)
frame@f9880000 = frame(4k)
frame@f9881000 = frame(4k)
frame@f9882000 = frame(4k)
frame@f9883000 = frame(4k)
frame@f9884000 = frame(4k)
frame@f9885000 = frame(4k)
frame@f9886000 = frame(4k)
frame@f9887000 = frame(4k)
frame@f9888000 = frame(4k)
frame@f9889000 = frame(4k)
frame@f988a000 = frame(4k)
frame@f988b000 = frame(4k)
frame@f988c000 = frame(4k)
frame@f988d000 = frame(4k)
frame@f988e000 = frame(4k)
frame@f988f000 = frame(4k)
frame@f9890000 = frame(4k)
frame@f9891000 = frame(4k)
frame@f9892000 = frame(4k)
frame@f9893000 = frame(4k)
frame@f9894000 = frame(4k)
frame@f9895000 = frame(4k)
frame@f9896000 = frame(4k)
frame@f9897000 = frame(4k)
frame@f9898000 = frame(4k)
frame@f9899000 = frame(4k)
frame@f989a000 = frame(4k)
frame@f989b000 = frame(4k)
frame@f989c000 = frame(4k)
frame@f989d000 = frame(4k)
frame@f989e000 = frame(4k)
frame@f989f000 = frame(4k)
frame@f98a0000 = frame(4k)
frame@f98a1000 = frame(4k)
frame@f98a2000 = frame(4k)
frame@f98a3000 = frame(4k)
frame@f98a4000 = frame(4k)
frame@f98a5000 = frame(4k)
frame@f98a6000 = frame(4k)
frame@f98a7000 = frame(4k)
frame@f98a8000 = frame(4k)
frame@f98a9000 = frame(4k)
frame@f98aa000 = frame(4k)
frame@f98ab000 = frame(4k)
frame@f98ac000 = frame(4k)
frame@f98ad000 = frame(4k)
frame@f98ae000 = frame(4k)
frame@f98af000 = frame(4k)
frame@f98b0000 = frame(4k)
frame@f98b1000 = frame(4k)
frame@f98b2000 = frame(4k)
frame@f98b3000 = frame(4k)
frame@f98b4000 = frame(4k)
frame@f98b5000 = frame(4k)
frame@f98b6000 = frame(4k)
frame@f98b7000 = frame(4k)
frame@f98b8000 = frame(4k)
frame@f98b9000 = frame(4k)
frame@f98ba000 = frame(4k)
frame@f98bb000 = frame(4k)
frame@f98bc000 = frame(4k)
frame@f98bd000 = frame(4k)
frame@f98be000 = frame(4k)
frame@f98bf000 = frame(4k)
frame@f98c0000 = frame(4k)
frame@f98c1000 = frame(4k)
frame@f98c2000 = frame(4k)
frame@f98c3000 = frame(4k)
frame@f98c4000 = frame(4k)
frame@f98c5000 = frame(4k)
frame@f98c6000 = frame(4k)
frame@f98c7000 = frame(4k)
frame@f98c8000 = frame(4k)
frame@f98c9000 = frame(4k)
frame@f98ca000 = frame(4k)
frame@f98cb000 = frame(4k)
frame@f98cc000 = frame(4k)
frame@f98cd000 = frame(4k)
frame@f98ce000 = frame(4k)
frame@f98cf000 = frame(4k)
frame@f98d0000 = frame(4k)
frame@f98d1000 = frame(4k)
frame@f98d2000 = frame(4k)
frame@f98d3000 = frame(4k)
frame@f98d4000 = frame(4k)
frame@f98d5000 = frame(4k)
frame@f98d6000 = frame(4k)
frame@f98d7000 = frame(4k)
frame@f98d8000 = frame(4k)
frame@f98d9000 = frame(4k)
frame@f98da000 = frame(4k)
frame@f98db000 = frame(4k)
frame@f98dc000 = frame(4k)
frame@f98dd000 = frame(4k)
frame@f98de000 = frame(4k)
frame@f98df000 = frame(4k)
frame@f98e0000 = frame(4k)
frame@f98e1000 = frame(4k)
frame@f98e2000 = frame(4k)
frame@f98e3000 = frame(4k)
frame@f98e4000 = frame(4k)
frame@f98e5000 = frame(4k)
frame@f98e6000 = frame(4k)
frame@f98e7000 = frame(4k)
frame@f98e8000 = frame(4k)
frame@f98e9000 = frame(4k)
frame@f98ea000 = frame(4k)
frame@f98eb000 = frame(4k)
frame@f98ec000 = frame(4k)
frame@f98ed000 = frame(4k)
frame@f98ee000 = frame(4k)
frame@f98ef000 = frame(4k)
frame@f98f0000 = frame(4k)
frame@f98f1000 = frame(4k)
frame@f98f2000 = frame(4k)
frame@f98f3000 = frame(4k)
frame@f98f4000 = frame(4k)
frame@f98f5000 = frame(4k)
frame@f98f6000 = frame(4k)
frame@f98f7000 = frame(4k)
frame@f98f8000 = frame(4k)
frame@f98f9000 = frame(4k)
frame@f98fa000 = frame(4k)
frame@f98fb000 = frame(4k)
frame@f98fc000 = frame(4k)
frame@f98fd000 = frame(4k)
frame@f98fe000 = frame(4k)
frame@f98ff000 = frame(4k)
frame@f9900000 = frame(4k)
frame@f9901000 = frame(4k)
frame@f9902000 = frame(4k)
frame@f9903000 = frame(4k)
frame@f9904000 = frame(4k)
frame@f9905000 = frame(4k)
frame@f9906000 = frame(4k)
frame@f9907000 = frame(4k)
frame@f9908000 = frame(4k)
frame@f9909000 = frame(4k)
frame@f990a000 = frame(4k)
frame@f990b000 = frame(4k)
frame@f990c000 = frame(4k)
frame@f990d000 = frame(4k)
frame@f990e000 = frame(4k)
frame@f990f000 = frame(4k)
frame@f9910000 = frame(4k)
frame@f9911000 = frame(4k)
frame@f9912000 = frame(4k)
frame@f9913000 = frame(4k)
frame@f9914000 = frame(4k)
frame@f9915000 = frame(4k)
frame@f9916000 = frame(4k)
frame@f9917000 = frame(4k)
frame@f9918000 = frame(4k)
frame@f9919000 = frame(4k)
frame@f991a000 = frame(4k)
frame@f991b000 = frame(4k)
frame@f991c000 = frame(4k)
frame@f991d000 = frame(4k)
frame@f991e000 = frame(4k)
frame@f991f000 = frame(4k)
frame@f9920000 = frame(4k)
frame@f9921000 = frame(4k)
frame@f9922000 = frame(4k)
frame@f9923000 = frame(4k)
frame@f9924000 = frame(4k)
frame@f9925000 = frame(4k)
frame@f9926000 = frame(4k)
frame@f9927000 = frame(4k)
frame@f9928000 = frame(4k)
frame@f9929000 = frame(4k)
frame@f992a000 = frame(4k)
frame@f992b000 = frame(4k)
frame@f992c000 = frame(4k)
frame@f992d000 = frame(4k)
frame@f992e000 = frame(4k)
frame@f992f000 = frame(4k)
frame@f9930000 = frame(4k)
frame@f9931000 = frame(4k)
frame@f9932000 = frame(4k)
frame@f9933000 = frame(4k)
frame@f9934000 = frame(4k)
frame@f9935000 = frame(4k)
frame@f9936000 = frame(4k)
frame@f9937000 = frame(4k)
frame@f9938000 = frame(4k)
frame@f9939000 = frame(4k)
frame@f993a000 = frame(4k)
frame@f993b000 = frame(4k)
frame@f993c000 = frame(4k)
frame@f993d000 = frame(4k)
frame@f993e000 = frame(4k)
frame@f993f000 = frame(4k)
frame@f9940000 = frame(4k)
frame@f9941000 = frame(4k)
frame@f9942000 = frame(4k)
frame@f9943000 = frame(4k)
frame@f9944000 = frame(4k)
frame@f9945000 = frame(4k)
frame@f9946000 = frame(4k)
frame@f9947000 = frame(4k)
frame@f9948000 = frame(4k)
frame@f9949000 = frame(4k)
frame@f994a000 = frame(4k)
frame@f994b000 = frame(4k)
frame@f994c000 = frame(4k)
frame@f994d000 = frame(4k)
frame@f994e000 = frame(4k)
frame@f994f000 = frame(4k)
frame@f9950000 = frame(4k)
frame@f9951000 = frame(4k)
frame@f9952000 = frame(4k)
frame@f9953000 = frame(4k)
frame@f9954000 = frame(4k)
frame@f9955000 = frame(4k)
frame@f9956000 = frame(4k)
frame@f9957000 = frame(4k)
frame@f9958000 = frame(4k)
frame@f9959000 = frame(4k)
frame@f995a000 = frame(4k)
frame@f995b000 = frame(4k)
frame@f995c000 = frame(4k)
frame@f995d000 = frame(4k)
frame@f995e000 = frame(4k)
frame@f995f000 = frame(4k)
frame@f9960000 = frame(4k)
frame@f9961000 = frame(4k)
frame@f9962000 = frame(4k)
frame@f9963000 = frame(4k)
frame@f9964000 = frame(4k)
frame@f9965000 = frame(4k)
frame@f9966000 = frame(4k)
frame@f9967000 = frame(4k)
frame@f9968000 = frame(4k)
frame@f9969000 = frame(4k)
frame@f996a000 = frame(4k)
frame@f996b000 = frame(4k)
frame@f996c000 = frame(4k)
frame@f996d000 = frame(4k)
frame@f996e000 = frame(4k)
frame@f996f000 = frame(4k)
frame@f9970000 = frame(4k)
frame@f9971000 = frame(4k)
frame@f9972000 = frame(4k)
frame@f9973000 = frame(4k)
frame@f9974000 = frame(4k)
frame@f9975000 = frame(4k)
frame@f9976000 = frame(4k)
frame@f9977000 = frame(4k)
frame@f9978000 = frame(4k)
frame@f9979000 = frame(4k)
frame@f997a000 = frame(4k)
frame@f997b000 = frame(4k)
frame@f997c000 = frame(4k)
frame@f997d000 = frame(4k)
frame@f997e000 = frame(4k)
frame@f997f000 = frame(4k)
frame@f9980000 = frame(4k)
frame@f9981000 = frame(4k)
frame@f9982000 = frame(4k)
frame@f9983000 = frame(4k)
frame@f9984000 = frame(4k)
frame@f9985000 = frame(4k)
frame@f9986000 = frame(4k)
frame@f9987000 = frame(4k)
frame@f9988000 = frame(4k)
frame@f9989000 = frame(4k)
frame@f998a000 = frame(4k)
frame@f998b000 = frame(4k)
frame@f998c000 = frame(4k)
frame@f998d000 = frame(4k)
frame@f998e000 = frame(4k)
frame@f998f000 = frame(4k)
frame@f9990000 = frame(4k)
frame@f9991000 = frame(4k)
frame@f9992000 = frame(4k)
frame@f9993000 = frame(4k)
frame@f9994000 = frame(4k)
frame@f9995000 = frame(4k)
frame@f9996000 = frame(4k)
frame@f9997000 = frame(4k)
frame@f9998000 = frame(4k)
frame@f9999000 = frame(4k)
frame@f999a000 = frame(4k)
frame@f999b000 = frame(4k)
frame@f999c000 = frame(4k)
frame@f999d000 = frame(4k)
frame@f999e000 = frame(4k)
frame@f999f000 = frame(4k)
frame@f99a0000 = frame(4k)
frame@f99a1000 = frame(4k)
frame@f99a2000 = frame(4k)
frame@f99a3000 = frame(4k)
frame@f99a4000 = frame(4k)
frame@f99a5000 = frame(4k)
frame@f99a6000 = frame(4k)
frame@f99a7000 = frame(4k)
frame@f99a8000 = frame(4k)
frame@f99a9000 = frame(4k)
frame@f99aa000 = frame(4k)
frame@f99ab000 = frame(4k)
frame@f99ac000 = frame(4k)
frame@f99ad000 = frame(4k)
frame@f99ae000 = frame(4k)
frame@f99af000 = frame(4k)
frame@f99b0000 = frame(4k)
frame@f99b1000 = frame(4k)
frame@f99b2000 = frame(4k)
frame@f99b3000 = frame(4k)
frame@f99b4000 = frame(4k)
frame@f99b5000 = frame(4k)
frame@f99b6000 = frame(4k)
frame@f99b7000 = frame(4k)
frame@f99b8000 = frame(4k)
frame@f99b9000 = frame(4k)
frame@f99ba000 = frame(4k)
frame@f99bb000 = frame(4k)
frame@f99bc000 = frame(4k)
frame@f99bd000 = frame(4k)
frame@f99be000 = frame(4k)
frame@f99bf000 = frame(4k)
frame@f99c0000 = frame(4k)
frame@f99c1000 = frame(4k)
frame@f99c2000 = frame(4k)
frame@f99c3000 = frame(4k)
frame@f99c4000 = frame(4k)
frame@f99c5000 = frame(4k)
frame@f99c6000 = frame(4k)
frame@f99c7000 = frame(4k)
frame@f99c8000 = frame(4k)
frame@f99c9000 = frame(4k)
frame@f99ca000 = frame(4k)
frame@f99cb000 = frame(4k)
frame@f99cc000 = frame(4k)
frame@f99cd000 = frame(4k)
frame@f99ce000 = frame(4k)
frame@f99cf000 = frame(4k)
frame@f99d0000 = frame(4k)
frame@f99d1000 = frame(4k)
frame@f99d2000 = frame(4k)
frame@f99d3000 = frame(4k)
frame@f99d4000 = frame(4k)
frame@f99d5000 = frame(4k)
frame@f99d6000 = frame(4k)
frame@f99d7000 = frame(4k)
frame@f99d8000 = frame(4k)
frame@f99d9000 = frame(4k)
frame@f99da000 = frame(4k)
frame@f99db000 = frame(4k)
frame@f99dc000 = frame(4k)
frame@f99dd000 = frame(4k)
frame@f99de000 = frame(4k)
frame@f99df000 = frame(4k)
frame@f99e0000 = frame(4k)
frame@f99e1000 = frame(4k)
frame@f99e2000 = frame(4k)
frame@f99e3000 = frame(4k)
frame@f99e4000 = frame(4k)
frame@f99e5000 = frame(4k)
frame@f99e6000 = frame(4k)
frame@f99e7000 = frame(4k)
frame@f99e8000 = frame(4k)
frame@f99e9000 = frame(4k)
frame@f99ea000 = frame(4k)
frame@f99eb000 = frame(4k)
frame@f99ec000 = frame(4k)
frame@f99ed000 = frame(4k)
frame@f99ee000 = frame(4k)
frame@f99ef000 = frame(4k)
frame@f99f0000 = frame(4k)
frame@f99f1000 = frame(4k)
frame@f99f2000 = frame(4k)
frame@f99f3000 = frame(4k)
frame@f99f4000 = frame(4k)
frame@f99f5000 = frame(4k)
frame@f99f6000 = frame(4k)
frame@f99f7000 = frame(4k)
frame@f99f8000 = frame(4k)
frame@f99f9000 = frame(4k)
frame@f99fa000 = frame(4k)
frame@f99fb000 = frame(4k)
frame@f99fc000 = frame(4k)
frame@f99fd000 = frame(4k)
frame@f99fe000 = frame(4k)
frame@f99ff000 = frame(4k)
frame@f9a00000 = frame(4k)
frame@f9a01000 = frame(4k)
frame@f9a02000 = frame(4k)
frame@f9a03000 = frame(4k)
frame@f9a04000 = frame(4k)
frame@f9a05000 = frame(4k)
frame@f9a06000 = frame(4k)
frame@f9a07000 = frame(4k)
frame@f9a08000 = frame(4k)
frame@f9a09000 = frame(4k)
frame@f9a0a000 = frame(4k)
frame@f9a0b000 = frame(4k)
frame@f9a0c000 = frame(4k)
frame@f9a0d000 = frame(4k)
frame@f9a0e000 = frame(4k)
frame@f9a0f000 = frame(4k)
frame@f9a10000 = frame(4k)
frame@f9a11000 = frame(4k)
frame@f9a12000 = frame(4k)
frame@f9a13000 = frame(4k)
frame@f9a14000 = frame(4k)
frame@f9a15000 = frame(4k)
frame@f9a16000 = frame(4k)
frame@f9a17000 = frame(4k)
frame@f9a18000 = frame(4k)
frame@f9a19000 = frame(4k)
frame@f9a1a000 = frame(4k)
frame@f9a1b000 = frame(4k)
frame@f9a1c000 = frame(4k)
frame@f9a1d000 = frame(4k)
frame@f9a1e000 = frame(4k)
frame@f9a1f000 = frame(4k)
frame@f9a20000 = frame(4k)
frame@f9a21000 = frame(4k)
frame@f9a22000 = frame(4k)
frame@f9a23000 = frame(4k)
frame@f9a24000 = frame(4k)
frame@f9a25000 = frame(4k)
frame@f9a26000 = frame(4k)
frame@f9a27000 = frame(4k)
frame@f9a28000 = frame(4k)
frame@f9a29000 = frame(4k)
frame@f9a2a000 = frame(4k)
frame@f9a2b000 = frame(4k)
frame@f9a2c000 = frame(4k)
frame@f9a2d000 = frame(4k)
frame@f9a2e000 = frame(4k)
frame@f9a2f000 = frame(4k)
frame@f9a30000 = frame(4k)
frame@f9a31000 = frame(4k)
frame@f9a32000 = frame(4k)
frame@f9a33000 = frame(4k)
frame@f9a34000 = frame(4k)
frame@f9a35000 = frame(4k)
frame@f9a36000 = frame(4k)
frame@f9a37000 = frame(4k)
frame@f9a38000 = frame(4k)
frame@f9a39000 = frame(4k)
frame@f9a3a000 = frame(4k)
frame@f9a3b000 = frame(4k)
frame@f9a3c000 = frame(4k)
frame@f9a3d000 = frame(4k)
frame@f9a3e000 = frame(4k)
frame@f9a3f000 = frame(4k)
frame@f9a40000 = frame(4k)
frame@f9a41000 = frame(4k)
frame@f9a42000 = frame(4k)
frame@f9a43000 = frame(4k)
frame@f9a44000 = frame(4k)
frame@f9a45000 = frame(4k)
frame@f9a46000 = frame(4k)
frame@f9a47000 = frame(4k)
frame@f9a48000 = frame(4k)
frame@f9a49000 = frame(4k)
frame@f9a4a000 = frame(4k)
frame@f9a4b000 = frame(4k)
frame@f9a4c000 = frame(4k)
frame@f9a4d000 = frame(4k)
frame@f9a4e000 = frame(4k)
frame@f9a4f000 = frame(4k)
frame@f9a50000 = frame(4k)
frame@f9a51000 = frame(4k)
frame@f9a52000 = frame(4k)
frame@f9a53000 = frame(4k)
frame@f9a54000 = frame(4k)
frame@f9a55000 = frame(4k)
frame@f9a56000 = frame(4k)
frame@f9a57000 = frame(4k)
frame@f9a58000 = frame(4k)
frame@f9a59000 = frame(4k)
frame@f9a5a000 = frame(4k)
frame@f9a5b000 = frame(4k)
frame@f9a5c000 = frame(4k)
frame@f9a5d000 = frame(4k)
frame@f9a5e000 = frame(4k)
frame@f9a5f000 = frame(4k)
frame@f9a60000 = frame(4k)
frame@f9a61000 = frame(4k)
frame@f9a62000 = frame(4k)
frame@f9a63000 = frame(4k)
frame@f9a64000 = frame(4k)
frame@f9a65000 = frame(4k)
frame@f9a66000 = frame(4k)
frame@f9a67000 = frame(4k)
frame@f9a68000 = frame(4k)
frame@f9a69000 = frame(4k)
frame@f9a6a000 = frame(4k)
frame@f9a6b000 = frame(4k)
frame@f9a6c000 = frame(4k)
frame@f9a6d000 = frame(4k)
frame@f9a6e000 = frame(4k)
frame@f9a6f000 = frame(4k)
frame@f9a70000 = frame(4k)
frame@f9a71000 = frame(4k)
frame@f9a72000 = frame(4k)
frame@f9a73000 = frame(4k)
frame@f9a74000 = frame(4k)
frame@f9a75000 = frame(4k)
frame@f9a76000 = frame(4k)
frame@f9a77000 = frame(4k)
frame@f9a78000 = frame(4k)
frame@f9a79000 = frame(4k)
frame@f9a7a000 = frame(4k)
frame@f9a7b000 = frame(4k)
frame@f9a7c000 = frame(4k)
frame@f9a7d000 = frame(4k)
frame@f9a7e000 = frame(4k)
frame@f9a7f000 = frame(4k)
frame@f9a80000 = frame(4k)
frame@f9a81000 = frame(4k)
frame@f9a82000 = frame(4k)
frame@f9a83000 = frame(4k)
frame@f9a84000 = frame(4k)
frame@f9a85000 = frame(4k)
frame@f9a86000 = frame(4k)
frame@f9a87000 = frame(4k)
frame@f9a88000 = frame(4k)
frame@f9a89000 = frame(4k)
frame@f9a8a000 = frame(4k)
frame@f9a8b000 = frame(4k)
frame@f9a8c000 = frame(4k)
frame@f9a8d000 = frame(4k)
frame@f9a8e000 = frame(4k)
frame@f9a8f000 = frame(4k)
frame@f9a90000 = frame(4k)
frame@f9a91000 = frame(4k)
frame@f9a92000 = frame(4k)
frame@f9a93000 = frame(4k)
frame@f9a94000 = frame(4k)
frame@f9a95000 = frame(4k)
frame@f9a96000 = frame(4k)
frame@f9a97000 = frame(4k)
frame@f9a98000 = frame(4k)
frame@f9a99000 = frame(4k)
frame@f9a9a000 = frame(4k)
frame@f9a9b000 = frame(4k)
frame@f9a9c000 = frame(4k)
frame@f9a9d000 = frame(4k)
frame@f9a9e000 = frame(4k)
frame@f9a9f000 = frame(4k)
frame@f9aa0000 = frame(4k)
frame@f9aa1000 = frame(4k)
frame@f9aa2000 = frame(4k)
frame@f9aa3000 = frame(4k)
frame@f9aa4000 = frame(4k)
frame@f9aa5000 = frame(4k)
frame@f9aa6000 = frame(4k)
frame@f9aa7000 = frame(4k)
frame@f9aa8000 = frame(4k)
frame@f9aa9000 = frame(4k)
frame@f9aaa000 = frame(4k)
frame@f9aab000 = frame(4k)
frame@f9aac000 = frame(4k)
frame@f9aad000 = frame(4k)
frame@f9aae000 = frame(4k)
frame@f9aaf000 = frame(4k)
frame@f9ab0000 = frame(4k)
frame@f9ab1000 = frame(4k)
frame@f9ab2000 = frame(4k)
frame@f9ab3000 = frame(4k)
frame@f9ab4000 = frame(4k)
frame@f9ab5000 = frame(4k)
frame@f9ab6000 = frame(4k)
frame@f9ab7000 = frame(4k)
frame@f9ab8000 = frame(4k)
frame@f9ab9000 = frame(4k)
frame@f9aba000 = frame(4k)
frame@f9abb000 = frame(4k)
frame@f9abc000 = frame(4k)
frame@f9abd000 = frame(4k)
frame@f9abe000 = frame(4k)
frame@f9abf000 = frame(4k)
frame@f9ac0000 = frame(4k)
frame@f9ac1000 = frame(4k)
frame@f9ac2000 = frame(4k)
frame@f9ac3000 = frame(4k)
frame@f9ac4000 = frame(4k)
frame@f9ac5000 = frame(4k)
frame@f9ac6000 = frame(4k)
frame@f9ac7000 = frame(4k)
frame@f9ac8000 = frame(4k)
frame@f9ac9000 = frame(4k)
frame@f9aca000 = frame(4k)
frame@f9acb000 = frame(4k)
frame@f9acc000 = frame(4k)
frame@f9acd000 = frame(4k)
frame@f9ace000 = frame(4k)
frame@f9acf000 = frame(4k)
frame@f9ad0000 = frame(4k)
frame@f9ad1000 = frame(4k)
frame@f9ad2000 = frame(4k)
frame@f9ad3000 = frame(4k)
frame@f9ad4000 = frame(4k)
frame@f9ad5000 = frame(4k)
frame@f9ad6000 = frame(4k)
frame@f9ad7000 = frame(4k)
frame@f9ad8000 = frame(4k)
frame@f9ad9000 = frame(4k)
frame@f9ada000 = frame(4k)
frame@f9adb000 = frame(4k)
frame@f9adc000 = frame(4k)
frame@f9add000 = frame(4k)
frame@f9ade000 = frame(4k)
frame@f9adf000 = frame(4k)
frame@f9ae0000 = frame(4k)
frame@f9ae1000 = frame(4k)
frame@f9ae2000 = frame(4k)
frame@f9ae3000 = frame(4k)
frame@f9ae4000 = frame(4k)
frame@f9ae5000 = frame(4k)
frame@f9ae6000 = frame(4k)
frame@f9ae7000 = frame(4k)
frame@f9ae8000 = frame(4k)
frame@f9ae9000 = frame(4k)
frame@f9aea000 = frame(4k)
frame@f9aeb000 = frame(4k)
frame@f9aec000 = frame(4k)
frame@f9aed000 = frame(4k)
frame@f9aee000 = frame(4k)
frame@f9aef000 = frame(4k)
frame@f9af0000 = frame(4k)
frame@f9af1000 = frame(4k)
frame@f9af2000 = frame(4k)
frame@f9af3000 = frame(4k)
frame@f9af4000 = frame(4k)
frame@f9af5000 = frame(4k)
frame@f9af6000 = frame(4k)
frame@f9af7000 = frame(4k)
frame@f9af8000 = frame(4k)
frame@f9af9000 = frame(4k)
frame@f9afa000 = frame(4k)
frame@f9afb000 = frame(4k)
frame@f9afc000 = frame(4k)
frame@f9afd000 = frame(4k)
frame@f9afe000 = frame(4k)
frame@f9aff000 = frame(4k)
frame@f9b00000 = frame(4k)
frame@f9b01000 = frame(4k)
frame@f9b02000 = frame(4k)
frame@f9b03000 = frame(4k)
frame@f9b04000 = frame(4k)
frame@f9b05000 = frame(4k)
frame@f9b06000 = frame(4k)
frame@f9b07000 = frame(4k)
frame@f9b08000 = frame(4k)
frame@f9b09000 = frame(4k)
frame@f9b0a000 = frame(4k)
frame@f9b0b000 = frame(4k)
frame@f9b0c000 = frame(4k)
frame@f9b0d000 = frame(4k)
frame@f9b0e000 = frame(4k)
frame@f9b0f000 = frame(4k)
frame@f9b10000 = frame(4k)
frame@f9b11000 = frame(4k)
frame@f9b12000 = frame(4k)
frame@f9b13000 = frame(4k)
frame@f9b14000 = frame(4k)
frame@f9b15000 = frame(4k)
frame@f9b16000 = frame(4k)
frame@f9b17000 = frame(4k)
frame@f9b18000 = frame(4k)
frame@f9b19000 = frame(4k)
frame@f9b1a000 = frame(4k)
frame@f9b1b000 = frame(4k)
frame@f9b1c000 = frame(4k)
frame@f9b1d000 = frame(4k)
frame@f9b1e000 = frame(4k)
frame@f9b1f000 = frame(4k)
frame@f9b20000 = frame(4k)
frame@f9b21000 = frame(4k)
frame@f9b22000 = frame(4k)
frame@f9b23000 = frame(4k)
frame@f9b24000 = frame(4k)
frame@f9b25000 = frame(4k)
frame@f9b26000 = frame(4k)
frame@f9b27000 = frame(4k)
frame@f9b28000 = frame(4k)
frame@f9b29000 = frame(4k)
frame@f9b2a000 = frame(4k)
frame@f9b2b000 = frame(4k)
frame@f9b2c000 = frame(4k)
frame@f9b2d000 = frame(4k)
frame@f9b2e000 = frame(4k)
frame@f9b2f000 = frame(4k)
frame@f9b30000 = frame(4k)
frame@f9b31000 = frame(4k)
frame@f9b32000 = frame(4k)
frame@f9b33000 = frame(4k)
frame@f9b34000 = frame(4k)
frame@f9b35000 = frame(4k)
frame@f9b36000 = frame(4k)
frame@f9b37000 = frame(4k)
frame@f9b38000 = frame(4k)
frame@f9b39000 = frame(4k)
frame@f9b3a000 = frame(4k)
frame@f9b3b000 = frame(4k)
frame@f9b3c000 = frame(4k)
frame@f9b3d000 = frame(4k)
frame@f9b3e000 = frame(4k)
frame@f9b3f000 = frame(4k)
frame@f9b40000 = frame(4k)
frame@f9b41000 = frame(4k)
frame@f9b42000 = frame(4k)
frame@f9b43000 = frame(4k)
frame@f9b44000 = frame(4k)
frame@f9b45000 = frame(4k)
frame@f9b46000 = frame(4k)
frame@f9b47000 = frame(4k)
frame@f9b48000 = frame(4k)
frame@f9b49000 = frame(4k)
frame@f9b4a000 = frame(4k)
frame@f9b4b000 = frame(4k)
frame@f9b4c000 = frame(4k)
frame@f9b4d000 = frame(4k)
frame@f9b4e000 = frame(4k)
frame@f9b4f000 = frame(4k)
frame@f9b50000 = frame(4k)
frame@f9b51000 = frame(4k)
frame@f9b52000 = frame(4k)
frame@f9b53000 = frame(4k)
frame@f9b54000 = frame(4k)
frame@f9b55000 = frame(4k)
frame@f9b56000 = frame(4k)
frame@f9b57000 = frame(4k)
frame@f9b58000 = frame(4k)
frame@f9b59000 = frame(4k)
frame@f9b5a000 = frame(4k)
frame@f9b5b000 = frame(4k)
frame@f9b5c000 = frame(4k)
frame@f9b5d000 = frame(4k)
frame@f9b5e000 = frame(4k)
frame@f9b5f000 = frame(4k)
frame@f9b60000 = frame(4k)
frame@f9b61000 = frame(4k)
frame@f9b62000 = frame(4k)
frame@f9b63000 = frame(4k)
frame@f9b64000 = frame(4k)
frame@f9b65000 = frame(4k)
frame@f9b66000 = frame(4k)
frame@f9b67000 = frame(4k)
frame@f9b68000 = frame(4k)
frame@f9b69000 = frame(4k)
frame@f9b6a000 = frame(4k)
frame@f9b6b000 = frame(4k)
frame@f9b6c000 = frame(4k)
frame@f9b6d000 = frame(4k)
frame@f9b6e000 = frame(4k)
frame@f9b6f000 = frame(4k)
frame@f9b70000 = frame(4k)
frame@f9b71000 = frame(4k)
frame@f9b72000 = frame(4k)
frame@f9b73000 = frame(4k)
frame@f9b74000 = frame(4k)
frame@f9b75000 = frame(4k)
frame@f9b76000 = frame(4k)
frame@f9b77000 = frame(4k)
frame@f9b78000 = frame(4k)
frame@f9b79000 = frame(4k)
frame@f9b7a000 = frame(4k)
frame@f9b7b000 = frame(4k)
frame@f9b7c000 = frame(4k)
frame@f9b7d000 = frame(4k)
frame@f9b7e000 = frame(4k)
frame@f9b7f000 = frame(4k)
frame@f9b80000 = frame(4k)
frame@f9b81000 = frame(4k)
frame@f9b82000 = frame(4k)
frame@f9b83000 = frame(4k)
frame@f9b84000 = frame(4k)
frame@f9b85000 = frame(4k)
frame@f9b86000 = frame(4k)
frame@f9b87000 = frame(4k)
frame@f9b88000 = frame(4k)
frame@f9b89000 = frame(4k)
frame@f9b8a000 = frame(4k)
frame@f9b8b000 = frame(4k)
frame@f9b8c000 = frame(4k)
frame@f9b8d000 = frame(4k)
frame@f9b8e000 = frame(4k)
frame@f9b8f000 = frame(4k)
frame@f9b90000 = frame(4k)
frame@f9b91000 = frame(4k)
frame@f9b92000 = frame(4k)
frame@f9b93000 = frame(4k)
frame@f9b94000 = frame(4k)
frame@f9b95000 = frame(4k)
frame@f9b96000 = frame(4k)
frame@f9b97000 = frame(4k)
frame@f9b98000 = frame(4k)
frame@f9b99000 = frame(4k)
frame@f9b9a000 = frame(4k)
frame@f9b9b000 = frame(4k)
frame@f9b9c000 = frame(4k)
frame@f9b9d000 = frame(4k)
frame@f9b9e000 = frame(4k)
frame@f9b9f000 = frame(4k)
frame@f9ba0000 = frame(4k)
frame@f9ba1000 = frame(4k)
frame@f9ba2000 = frame(4k)
frame@f9ba3000 = frame(4k)
frame@f9ba4000 = frame(4k)
frame@f9ba5000 = frame(4k)
frame@f9ba6000 = frame(4k)
frame@f9ba7000 = frame(4k)
frame@f9ba8000 = frame(4k)
frame@f9ba9000 = frame(4k)
frame@f9baa000 = frame(4k)
frame@f9bab000 = frame(4k)
frame@f9bac000 = frame(4k)
frame@f9bad000 = frame(4k)
frame@f9bae000 = frame(4k)
frame@f9baf000 = frame(4k)
frame@f9bb0000 = frame(4k)
frame@f9bb1000 = frame(4k)
frame@f9bb2000 = frame(4k)
frame@f9bb3000 = frame(4k)
frame@f9bb4000 = frame(4k)
frame@f9bb5000 = frame(4k)
frame@f9bb6000 = frame(4k)
frame@f9bb7000 = frame(4k)
frame@f9bb8000 = frame(4k)
frame@f9bb9000 = frame(4k)
frame@f9bba000 = frame(4k)
frame@f9bbb000 = frame(4k)
frame@f9bbc000 = frame(4k)
frame@f9bbd000 = frame(4k)
frame@f9bbe000 = frame(4k)
frame@f9bbf000 = frame(4k)
frame@f9bc0000 = frame(4k)
frame@f9bc1000 = frame(4k)
frame@f9bc2000 = frame(4k)
frame@f9bc3000 = frame(4k)
frame@f9bc4000 = frame(4k)
frame@f9bc5000 = frame(4k)
frame@f9bc6000 = frame(4k)
frame@f9bc7000 = frame(4k)
frame@f9bc8000 = frame(4k)
frame@f9bc9000 = frame(4k)
frame@f9bca000 = frame(4k)
frame@f9bcb000 = frame(4k)
frame@f9bcc000 = frame(4k)
frame@f9bcd000 = frame(4k)
frame@f9bce000 = frame(4k)
frame@f9bcf000 = frame(4k)
frame@f9bd0000 = frame(4k)
frame@f9bd1000 = frame(4k)
frame@f9bd2000 = frame(4k)
frame@f9bd3000 = frame(4k)
frame@f9bd4000 = frame(4k)
frame@f9bd5000 = frame(4k)
frame@f9bd6000 = frame(4k)
frame@f9bd7000 = frame(4k)
frame@f9bd8000 = frame(4k)
frame@f9bd9000 = frame(4k)
frame@f9bda000 = frame(4k)
frame@f9bdb000 = frame(4k)
frame@f9bdc000 = frame(4k)
frame@f9bdd000 = frame(4k)
frame@f9bde000 = frame(4k)
frame@f9bdf000 = frame(4k)
frame@f9be0000 = frame(4k)
frame@f9be1000 = frame(4k)
frame@f9be2000 = frame(4k)
frame@f9be3000 = frame(4k)
frame@f9be4000 = frame(4k)
frame@f9be5000 = frame(4k)
frame@f9be6000 = frame(4k)
frame@f9be7000 = frame(4k)
frame@f9be8000 = frame(4k)
frame@f9be9000 = frame(4k)
frame@f9bea000 = frame(4k)
frame@f9beb000 = frame(4k)
frame@f9bec000 = frame(4k)
frame@f9bed000 = frame(4k)
frame@f9bee000 = frame(4k)
frame@f9bef000 = frame(4k)
frame@f9bf0000 = frame(4k)
frame@f9bf1000 = frame(4k)
frame@f9bf2000 = frame(4k)
frame@f9bf3000 = frame(4k)
frame@f9bf4000 = frame(4k)
frame@f9bf5000 = frame(4k)
frame@f9bf6000 = frame(4k)
frame@f9bf7000 = frame(4k)
frame@f9bf8000 = frame(4k)
frame@f9bf9000 = frame(4k)
frame@f9bfa000 = frame(4k)
frame@f9bfb000 = frame(4k)
frame@f9bfc000 = frame(4k)
frame@f9bfd000 = frame(4k)
frame@f9bfe000 = frame(4k)
frame@f9bff000 = frame(4k)
frame@f9c00000 = frame(4k)
frame@f9c01000 = frame(4k)
frame@f9c02000 = frame(4k)
frame@f9c03000 = frame(4k)
frame@f9c04000 = frame(4k)
frame@f9c05000 = frame(4k)
frame@f9c06000 = frame(4k)
frame@f9c07000 = frame(4k)
frame@f9c08000 = frame(4k)
frame@f9c09000 = frame(4k)
frame@f9c0a000 = frame(4k)
frame@f9c0b000 = frame(4k)
frame@f9c0c000 = frame(4k)
frame@f9c0d000 = frame(4k)
frame@f9c0e000 = frame(4k)
frame@f9c0f000 = frame(4k)
frame@f9c10000 = frame(4k)
frame@f9c11000 = frame(4k)
frame@f9c12000 = frame(4k)
frame@f9c13000 = frame(4k)
frame@f9c14000 = frame(4k)
frame@f9c15000 = frame(4k)
frame@f9c16000 = frame(4k)
frame@f9c17000 = frame(4k)
frame@f9c18000 = frame(4k)
frame@f9c19000 = frame(4k)
frame@f9c1a000 = frame(4k)
frame@f9c1b000 = frame(4k)
frame@f9c1c000 = frame(4k)
frame@f9c1d000 = frame(4k)
frame@f9c1e000 = frame(4k)
frame@f9c1f000 = frame(4k)
frame@f9c20000 = frame(4k)
frame@f9c21000 = frame(4k)
frame@f9c22000 = frame(4k)
frame@f9c23000 = frame(4k)
frame@f9c24000 = frame(4k)
frame@f9c25000 = frame(4k)
frame@f9c26000 = frame(4k)
frame@f9c27000 = frame(4k)
frame@f9c28000 = frame(4k)
frame@f9c29000 = frame(4k)
frame@f9c2a000 = frame(4k)
frame@f9c2b000 = frame(4k)
frame@f9c2c000 = frame(4k)
frame@f9c2d000 = frame(4k)
frame@f9c2e000 = frame(4k)
frame@f9c2f000 = frame(4k)
frame@f9c30000 = frame(4k)
frame@f9c31000 = frame(4k)
frame@f9c32000 = frame(4k)
frame@f9c33000 = frame(4k)
frame@f9c34000 = frame(4k)
frame@f9c35000 = frame(4k)
frame@f9c36000 = frame(4k)
frame@f9c37000 = frame(4k)
frame@f9c38000 = frame(4k)
frame@f9c39000 = frame(4k)
frame@f9c3a000 = frame(4k)
frame@f9c3b000 = frame(4k)
frame@f9c3c000 = frame(4k)
frame@f9c3d000 = frame(4k)
frame@f9c3e000 = frame(4k)
frame@f9c3f000 = frame(4k)
frame@f9c40000 = frame(4k)
frame@f9c41000 = frame(4k)
frame@f9c42000 = frame(4k)
frame@f9c43000 = frame(4k)
frame@f9c44000 = frame(4k)
frame@f9c45000 = frame(4k)
frame@f9c46000 = frame(4k)
frame@f9c47000 = frame(4k)
frame@f9c48000 = frame(4k)
frame@f9c49000 = frame(4k)
frame@f9c4a000 = frame(4k)
frame@f9c4b000 = frame(4k)
frame@f9c4c000 = frame(4k)
frame@f9c4d000 = frame(4k)
frame@f9c4e000 = frame(4k)
frame@f9c4f000 = frame(4k)
frame@f9c50000 = frame(4k)
frame@f9c51000 = frame(4k)
frame@f9c52000 = frame(4k)
frame@f9c53000 = frame(4k)
frame@f9c54000 = frame(4k)
frame@f9c55000 = frame(4k)
frame@f9c56000 = frame(4k)
frame@f9c57000 = frame(4k)
frame@f9c58000 = frame(4k)
frame@f9c59000 = frame(4k)
frame@f9c5a000 = frame(4k)
frame@f9c5b000 = frame(4k)
frame@f9c5c000 = frame(4k)
frame@f9c5d000 = frame(4k)
frame@f9c5e000 = frame(4k)
frame@f9c5f000 = frame(4k)
frame@f9c60000 = frame(4k)
frame@f9c61000 = frame(4k)
frame@f9c62000 = frame(4k)
frame@f9c63000 = frame(4k)
frame@f9c64000 = frame(4k)
frame@f9c65000 = frame(4k)
frame@f9c66000 = frame(4k)
frame@f9c67000 = frame(4k)
frame@f9c68000 = frame(4k)
frame@f9c69000 = frame(4k)
frame@f9c6a000 = frame(4k)
frame@f9c6b000 = frame(4k)
frame@f9c6c000 = frame(4k)
frame@f9c6d000 = frame(4k)
frame@f9c6e000 = frame(4k)
frame@f9c6f000 = frame(4k)
frame@f9c70000 = frame(4k)
frame@f9c71000 = frame(4k)
frame@f9c72000 = frame(4k)
frame@f9c73000 = frame(4k)
frame@f9c74000 = frame(4k)
frame@f9c75000 = frame(4k)
frame@f9c76000 = frame(4k)
frame@f9c77000 = frame(4k)
frame@f9c78000 = frame(4k)
frame@f9c79000 = frame(4k)
frame@f9c7a000 = frame(4k)
frame@f9c7b000 = frame(4k)
frame@f9c7c000 = frame(4k)
frame@f9c7d000 = frame(4k)
frame@f9c7e000 = frame(4k)
frame@f9c7f000 = frame(4k)
frame@f9c80000 = frame(4k)
frame@f9c81000 = frame(4k)
frame@f9c82000 = frame(4k)
frame@f9c83000 = frame(4k)
frame@f9c84000 = frame(4k)
frame@f9c85000 = frame(4k)
frame@f9c86000 = frame(4k)
frame@f9c87000 = frame(4k)
frame@f9c88000 = frame(4k)
frame@f9c89000 = frame(4k)
frame@f9c8a000 = frame(4k)
frame@f9c8b000 = frame(4k)
frame@f9c8c000 = frame(4k)
frame@f9c8d000 = frame(4k)
frame@f9c8e000 = frame(4k)
frame@f9c8f000 = frame(4k)
frame@f9c90000 = frame(4k)
frame@f9c91000 = frame(4k)
frame@f9c92000 = frame(4k)
frame@f9c93000 = frame(4k)
frame@f9c94000 = frame(4k)
frame@f9c95000 = frame(4k)
frame@f9c96000 = frame(4k)
frame@f9c97000 = frame(4k)
frame@f9c98000 = frame(4k)
frame@f9c99000 = frame(4k)
frame@f9c9a000 = frame(4k)
frame@f9c9b000 = frame(4k)
frame@f9c9c000 = frame(4k)
frame@f9c9d000 = frame(4k)
frame@f9c9e000 = frame(4k)
frame@f9c9f000 = frame(4k)
frame@f9ca0000 = frame(4k)
frame@f9ca1000 = frame(4k)
frame@f9ca2000 = frame(4k)
frame@f9ca3000 = frame(4k)
frame@f9ca4000 = frame(4k)
frame@f9ca5000 = frame(4k)
frame@f9ca6000 = frame(4k)
frame@f9ca7000 = frame(4k)
frame@f9ca8000 = frame(4k)
frame@f9ca9000 = frame(4k)
frame@f9caa000 = frame(4k)
frame@f9cab000 = frame(4k)
frame@f9cac000 = frame(4k)
frame@f9cad000 = frame(4k)
frame@f9cae000 = frame(4k)
frame@f9caf000 = frame(4k)
frame@f9cb0000 = frame(4k)
frame@f9cb1000 = frame(4k)
frame@f9cb2000 = frame(4k)
frame@f9cb3000 = frame(4k)
frame@f9cb4000 = frame(4k)
frame@f9cb5000 = frame(4k)
frame@f9cb6000 = frame(4k)
frame@f9cb7000 = frame(4k)
frame@f9cb8000 = frame(4k)
frame@f9cb9000 = frame(4k)
frame@f9cba000 = frame(4k)
frame@f9cbb000 = frame(4k)
frame@f9cbc000 = frame(4k)
frame@f9cbd000 = frame(4k)
frame@f9cbe000 = frame(4k)
frame@f9cbf000 = frame(4k)
frame@f9cc0000 = frame(4k)
frame@f9cc1000 = frame(4k)
frame@f9cc2000 = frame(4k)
frame@f9cc3000 = frame(4k)
frame@f9cc4000 = frame(4k)
frame@f9cc5000 = frame(4k)
frame@f9cc6000 = frame(4k)
frame@f9cc7000 = frame(4k)
frame@f9cc8000 = frame(4k)
frame@f9cc9000 = frame(4k)
frame@f9cca000 = frame(4k)
frame@f9ccb000 = frame(4k)
frame@f9ccc000 = frame(4k)
frame@f9ccd000 = frame(4k)
frame@f9cce000 = frame(4k)
frame@f9ccf000 = frame(4k)
frame@f9cd0000 = frame(4k)
frame@f9cd1000 = frame(4k)
frame@f9cd2000 = frame(4k)
frame@f9cd3000 = frame(4k)
frame@f9cd4000 = frame(4k)
frame@f9cd5000 = frame(4k)
frame@f9cd6000 = frame(4k)
frame@f9cd7000 = frame(4k)
frame@f9cd8000 = frame(4k)
frame@f9cd9000 = frame(4k)
frame@f9cda000 = frame(4k)
frame@f9cdb000 = frame(4k)
frame@f9cdc000 = frame(4k)
frame@f9cdd000 = frame(4k)
frame@f9cde000 = frame(4k)
frame@f9cdf000 = frame(4k)
frame@f9ce0000 = frame(4k)
frame@f9ce1000 = frame(4k)
frame@f9ce2000 = frame(4k)
frame@f9ce3000 = frame(4k)
frame@f9ce4000 = frame(4k)
frame@f9ce5000 = frame(4k)
frame@f9ce6000 = frame(4k)
frame@f9ce7000 = frame(4k)
frame@f9ce8000 = frame(4k)
frame@f9ce9000 = frame(4k)
frame@f9cea000 = frame(4k)
frame@f9ceb000 = frame(4k)
frame@f9cec000 = frame(4k)
frame@f9ced000 = frame(4k)
frame@f9cee000 = frame(4k)
frame@f9cef000 = frame(4k)
frame@f9cf0000 = frame(4k)
frame@f9cf1000 = frame(4k)
frame@f9cf2000 = frame(4k)
frame@f9cf3000 = frame(4k)
frame@f9cf4000 = frame(4k)
frame@f9cf5000 = frame(4k)
frame@f9cf6000 = frame(4k)
frame@f9cf7000 = frame(4k)
frame@f9cf8000 = frame(4k)
frame@f9cf9000 = frame(4k)
frame@f9cfa000 = frame(4k)
frame@f9cfb000 = frame(4k)
frame@f9cfc000 = frame(4k)
frame@f9cfd000 = frame(4k)
frame@f9cfe000 = frame(4k)
frame@f9cff000 = frame(4k)
frame@f9dc2000 = frame(4k)
frame@f9dc3000 = frame(4k)
frame@f9dc4000 = frame(4k)
frame@f9dc5000 = frame(4k)
frame@f9dc6000 = frame(4k)
frame@f9dc7000 = frame(4k)
frame@f9dc8000 = frame(4k)
frame@f9dc9000 = frame(4k)
frame@f9dca000 = frame(4k)
frame@f9dcb000 = frame(4k)
frame@f9dcc000 = frame(4k)
frame@f9dcd000 = frame(4k)
frame@f9dce000 = frame(4k)
frame@f9dcf000 = frame(4k)
frame@f9dd0000 = frame(4k)
frame@f9dd1000 = frame(4k)
frame@f9dd2000 = frame(4k)
frame@f9dd3000 = frame(4k)
frame@f9dd4000 = frame(4k)
frame@f9dd5000 = frame(4k)
frame@f9dd6000 = frame(4k)
frame@f9dd7000 = frame(4k)
frame@f9dd8000 = frame(4k)
frame@f9dd9000 = frame(4k)
frame@f9dda000 = frame(4k)
frame@f9ddb000 = frame(4k)
frame@f9ddc000 = frame(4k)
frame@f9ddd000 = frame(4k)
frame@f9dde000 = frame(4k)
frame@f9ddf000 = frame(4k)
frame@f9de0000 = frame(4k)
frame@f9de1000 = frame(4k)
frame@f9de2000 = frame(4k)
frame@f9de3000 = frame(4k)
frame@f9de4000 = frame(4k)
frame@f9de5000 = frame(4k)
frame@f9de6000 = frame(4k)
frame@f9de7000 = frame(4k)
frame@f9de8000 = frame(4k)
frame@f9de9000 = frame(4k)
frame@f9dea000 = frame(4k)
frame@f9deb000 = frame(4k)
frame@f9dec000 = frame(4k)
frame@f9ded000 = frame(4k)
frame@f9dee000 = frame(4k)
frame@f9def000 = frame(4k)
frame@f9df0000 = frame(4k)
frame@f9df1000 = frame(4k)
frame@f9df2000 = frame(4k)
frame@f9df3000 = frame(4k)
frame@f9df4000 = frame(4k)
frame@f9df5000 = frame(4k)
frame@f9df6000 = frame(4k)
frame@f9df7000 = frame(4k)
frame@f9df8000 = frame(4k)
frame@f9df9000 = frame(4k)
frame@f9dfa000 = frame(4k)
frame@f9dfb000 = frame(4k)
frame@f9dfc000 = frame(4k)
frame@f9dfd000 = frame(4k)
frame@f9dfe000 = frame(4k)
frame@f9dff000 = frame(4k)
pt@f6df3000 = pt
pt@f6df4000 = pt
pt@f6df5000 = pt
pt@f6df6000 = pt
pt@f6df7000 = pt
pt@f6df8000 = pt
pt@f6df9000 = pt
pt@f6dfa000 = pt
pt@f6dfb000 = pt
pt@f6dfc000 = pt
pt@f6dfd000 = pt
pt@f6dff000 = pt
pd@f6c7c000 = pd
pd@f6c7d000 = pd
pd@f6c7e000 = pd
pd@f6c7f000 = pd
irqhandler@0 = irq
irqhandler@19 = irq
irqhandler@1a = irq
irqhandler@1b = irq
irqhandler@1c = irq
asid_pool@e0130000 = asid_pool
asid_pool@e0132000 = asid_pool
asid_pool@e182f000 = asid_pool
iospace@c8 = io_device
iospace@100 = io_device
iospace@101 = io_device
iospace@2000 = io_device

caps

tcb@fffeed00{
  0: cnode@f6bf4000
  1: pd@f6c7f000
  2: tcb@fffeed00(reply)
  4: frame@f6cff000
}
tcb@fffee900{
  0: cnode@f6bf0000
  1: pd@f6c7e000
  2: tcb@fffee900(reply)
  4: frame@f6cf1000
}
tcb@fffee500{
  0: cnode@f6bcc000
  1: pd@f6c7c000
  2: tcb@fffee500(reply)
  4: frame@f729d000
}
cnode@f6bf4000{
  1: tcb@fffeed00
  2: cnode@f6bf4000
  3: pd@f6c7f000
  6: asid_pool@e0130000
  11: untyped@e0131000@12
  12: irqhandler@0
  13: ioports (ports: [64..67])
  14: aep@fffeffd0 (badge: 0x4, W )
  15: aep@fffeffe0 (badge: 0x10, W )
}
cnode@f6bf0000{
  1: tcb@fffee900
  2: cnode@f6bf0000 
  3: pd@f6c7e000
  6: asid_pool@e0132000
  11: pd@f6c7d000
  12: untyped@e0133000@12
  13: untyped@e0134000@12
  14: untyped@e0135000@12
  15: untyped@e0136000@12
  16: untyped@e0137000@12
  17: untyped@e0138000@12
  18: untyped@e0139000@12
  19: untyped@e013a000@12
  20: untyped@e013b000@12
  21: untyped@e013c000@12
  22: untyped@e013d000@12
  23: untyped@e013e000@12
  24: untyped@e013f000@12
  25: untyped@e0030000@12
  26: untyped@e0031000@12
  27: untyped@e0032000@12
  28: untyped@e0033000@12
  29: untyped@e0034000@12
  30: untyped@e0035000@12
  31: untyped@e0036000@12
  32: untyped@e0037000@12
  33: untyped@e0038000@12
  34: untyped@e0039000@12
  35: untyped@e003a000@12
  36: untyped@e003b000@12
  37: untyped@e003c000@12
  38: untyped@e003d000@12
  39: untyped@e003e000@12
  40: untyped@e003f000@12
  41: untyped@e0c40000@12
  42: untyped@e0c41000@12
  43: untyped@e0c42000@12
  44: untyped@e0c43000@12
  45: untyped@e0c44000@12
  46: untyped@e0c45000@12
  47: untyped@e0c46000@12
  48: untyped@e0c47000@12
  49: untyped@e0028000@12
  50: untyped@e0029000@12
  51: untyped@e002a000@12
  52: untyped@e002b000@12
  53: untyped@e002c000@12
  54: untyped@e002d000@12
  55: untyped@e002e000@12
  56: untyped@e002f000@12
  57: untyped@e0090000@12
  58: untyped@e0091000@12
  59: untyped@e0092000@12
  60: untyped@e0093000@12
  61: untyped@e182e000@12
  62: untyped@f7300000@20
  63: untyped@f7400000@20
  64: untyped@f7500000@20
  65: untyped@f7600000@20
  66: untyped@f7700000@20
  67: untyped@f7800000@20
  68: untyped@f7900000@20
  69: untyped@f7a00000@20
  70: untyped@f7b00000@20
  71: untyped@f7c00000@20
  72: untyped@f7d00000@20
  73: untyped@f7e00000@20
  74: untyped@f7f00000@20
  75: untyped@e4000000@20
  76: untyped@e4100000@20
  77: untyped@e4200000@20
  78: untyped@e4300000@20
  79: untyped@e4400000@20
  80: untyped@e4500000@20
  81: untyped@e4600000@20
  82: untyped@e4700000@20
  83: untyped@e4800000@20
  84: untyped@e4900000@20
  85: untyped@e4a00000@20
  86: untyped@e4b00000@20
  87: untyped@e4c00000@20
  88: untyped@e4d00000@20
  89: untyped@e4e00000@20
  90: untyped@e4f00000@20
  91: untyped@e5000000@20
  92: untyped@e5100000@20
  93: untyped@e5200000@20
  94: untyped@e5300000@20
  95: untyped@e5400000@20
  96: untyped@e5500000@20
  97: untyped@e5600000@20
  98: untyped@e5700000@20
  99: untyped@e5800000@20
  100: untyped@e5900000@20
  101: untyped@e5a00000@20
  102: untyped@e5b00000@20
  103: untyped@e5c00000@20
  104: untyped@e5d00000@20
  105: untyped@e5e00000@20
  106: untyped@e5f00000@20
  107: untyped@e6000000@20
  108: untyped@e6100000@20
  109: untyped@e6200000@20
  110: untyped@e6300000@20
  111: untyped@e6400000@20
  112: untyped@e6500000@20
  113: untyped@e6600000@20
  114: untyped@e6700000@20
  115: untyped@e6800000@20
  116: untyped@e6900000@20
  117: untyped@e6a00000@20
  118: untyped@e6b00000@20
  119: untyped@e6c00000@20
  120: untyped@e6d00000@20
  121: untyped@e6e00000@20
  122: untyped@e6f00000@20
  123: untyped@e7000000@20
  124: untyped@e7100000@20
  125: untyped@e7200000@20
  126: untyped@e7300000@20
  127: untyped@e7400000@20
  128: untyped@e7500000@20
  129: untyped@e7600000@20
  130: untyped@e7700000@20
  131: untyped@e7800000@20
  132: untyped@e7900000@20
  133: untyped@e7a00000@20
  134: untyped@e7b00000@20
  135: untyped@e7c00000@20
  136: untyped@e7d00000@20
  137: untyped@e7e00000@20
  138: untyped@e7f00000@20
  139: untyped@f8000000@20
  140: untyped@f8100000@20
  141: untyped@f8200000@20
  142: untyped@f8300000@20
  143: untyped@f8400000@20
  144: untyped@f8500000@20
  145: untyped@f8600000@20
  146: untyped@f8700000@20
  147: untyped@f8800000@20
  148: untyped@f8900000@20
  149: untyped@f8a00000@20
  150: untyped@f8b00000@20
  151: untyped@f8c00000@20
  152: untyped@f8d00000@20
  153: untyped@f8e00000@20
  154: untyped@f8f00000@20
  155: untyped@f9000000@20
  156: untyped@f9100000@20
  157: untyped@f9200000@20
  158: untyped@f9300000@20
  159: untyped@f9400000@20
  160: untyped@f9500000@20
  161: untyped@f9600000@20
  162: untyped@f9700000@20
  163: irqhandler@19
  164: frame@d0200000
  165: frame@d0201000
  166: frame@d0202000
  167: frame@d0203000
  168: frame@d0204000
  169: frame@d0205000
  170: frame@d0206000
  171: frame@d0207000
  172: frame@d0208000
  173: frame@d0209000
  174: frame@d020a000
  175: frame@d020b000
  176: frame@d020c000
  177: frame@d020d000
  178: frame@d020e000
  179: frame@d020f000
  180: frame@d0210000
  181: frame@d0211000
  182: frame@d0212000
  183: frame@d0213000
  184: frame@d0214000
  185: frame@d0215000
  186: frame@d0216000
  187: frame@d0217000
  188: frame@d0218000
  189: frame@d0219000
  190: frame@d021a000
  191: frame@d021b000
  192: frame@d021c000
  193: frame@d021d000
  194: frame@d021e000
  195: frame@d021f000
  196: frame@d0220000
  197: frame@d0221000
  198: frame@d0222000
  199: frame@d0223000
  200: frame@d0224000
  201: frame@d0225000
  202: frame@d0226000
  203: frame@d0227000
  204: frame@d0228000
  205: frame@d0229000
  206: frame@d022a000
  207: frame@d022b000
  208: frame@d022c000
  209: frame@d022d000
  210: frame@d022e000
  211: frame@d022f000
  212: frame@d0230000
  213: frame@d0231000
  214: frame@d0232000
  215: frame@d0233000
  216: frame@d0234000
  217: frame@d0235000
  218: frame@d0236000
  219: frame@d0237000
  220: frame@d0238000
  221: frame@d0239000
  222: frame@d023a000
  223: frame@d023b000
  224: frame@d023c000
  225: frame@d023d000
  226: frame@d023e000
  227: frame@d023f000
  228: iospace@100
  229: irqhandler@1a
  230: frame@d0240000
  231: frame@d0241000
  232: frame@d0242000
  233: frame@d0243000
  234: frame@d0244000
  235: frame@d0245000
  236: frame@d0246000
  237: frame@d0247000
  238: frame@d0248000
  239: frame@d0249000
  240: frame@d024a000
  241: frame@d024b000
  242: frame@d024c000
  243: frame@d024d000
  244: frame@d024e000
  245: frame@d024f000
  246: frame@d0250000
  247: frame@d0251000
  248: frame@d0252000
  249: frame@d0253000
  250: frame@d0254000
  251: frame@d0255000
  252: frame@d0256000
  253: frame@d0257000
  254: frame@d0258000
  255: frame@d0259000
  256: frame@d025a000
  257: frame@d025b000
  258: frame@d025c000
  259: frame@d025d000
  260: frame@d025e000
  261: frame@d025f000
  262: frame@d0260000
  263: frame@d0261000
  264: frame@d0262000
  265: frame@d0263000
  266: frame@d0264000
  267: frame@d0265000
  268: frame@d0266000
  269: frame@d0267000
  270: frame@d0268000
  271: frame@d0269000
  272: frame@d026a000
  273: frame@d026b000
  274: frame@d026c000
  275: frame@d026d000
  276: frame@d026e000
  277: frame@d026f000
  278: frame@d0270000
  279: frame@d0271000
  280: frame@d0272000
  281: frame@d0273000
  282: frame@d0274000
  283: frame@d0275000
  284: frame@d0276000
  285: frame@d0277000
  286: frame@d0278000
  287: frame@d0279000
  288: frame@d027a000
  289: frame@d027b000
  290: frame@d027c000
  291: frame@d027d000
  292: frame@d027e000
  293: frame@d027f000
  294: iospace@101
  295: irqhandler@1c
  296: frame@d0300000
  297: frame@d0301000
  298: frame@d0302000
  299: frame@d0303000
  300: iospace@2000
  301: ioports (ports: [3320..3327])
  302: ep@e001cff0 (  R)
  303: aep@fffeffe0 (badge: 0x0,  R)
}
cnode@f6bc8000{
  1: tcb@fffee500
  2: cnode@f6bcc000
  3: pd@f6c7c000
  6: asid_pool@e182f000
  11: untyped@e0c48000@12
  12: untyped@e0c49000@12
  13: untyped@e012e000@12
  14: untyped@e012f000@12
  15: untyped@e0026000@12
  16: untyped@e0027000@12
  17: untyped@e009c000@12
  18: untyped@e009d000@12
  19: untyped@e182d000@12
  20: untyped@e009e000@12
  21: untyped@e0022000@12
  22: untyped@e0021000@12
  23: untyped@e0020000@12
  24: untyped@e001f000@12
  25: untyped@e001e000@12
  26: untyped@e001d000@12
  27: untyped@f9e00000@20
  28: untyped@f9f00000@20
  29: untyped@fa000000@20
  30: untyped@fa100000@20
  31: untyped@fa200000@20
  32: untyped@fa300000@20
  33: untyped@fa400000@20
  34: untyped@fa500000@20
  35: untyped@fa600000@20
  36: untyped@fa700000@20
  37: untyped@fa800000@20
  38: untyped@fa900000@20
  39: untyped@faa00000@20
  40: untyped@fab00000@20
  41: untyped@fac00000@20
  42: untyped@fad00000@20
  43: untyped@fae00000@20
  44: untyped@faf00000@20
  45: untyped@fb000000@20
  46: untyped@fb100000@20
  47: untyped@fb200000@20
  48: untyped@fb300000@20
  49: untyped@fb400000@20
  50: untyped@fb500000@20
  51: untyped@fb600000@20
  52: untyped@fb700000@20
  53: untyped@fb800000@20
  54: untyped@fb900000@20
  55: untyped@fba00000@20
  56: untyped@fbb00000@20
  57: untyped@fbc00000@20
  58: untyped@fbd00000@20
  59: untyped@fbe00000@20
  60: untyped@fbf00000@20
  61: untyped@e2000000@20
  62: untyped@e2100000@20
  63: untyped@e2200000@20
  64: untyped@e2300000@20
  65: untyped@e2400000@20
  66: untyped@e2500000@20
  67: untyped@e2600000@20
  68: untyped@e2700000@20
  69: untyped@e2800000@20
  70: untyped@e2900000@20
  71: untyped@e2a00000@20
  72: untyped@e2b00000@20
  73: untyped@e2c00000@20
  74: untyped@e2d00000@20
  75: untyped@e2e00000@20
  76: untyped@e2f00000@20
  77: untyped@e3000000@20
  78: untyped@e3100000@20
  79: untyped@e3200000@20
  80: untyped@e3300000@20
  81: untyped@e3400000@20
  82: untyped@e3500000@20
  83: untyped@e3600000@20
  84: untyped@e3700000@20
  85: untyped@e3800000@20
  86: untyped@e3900000@20
  87: untyped@e3a00000@20
  88: untyped@e3b00000@20
  89: untyped@e3c00000@20
  90: untyped@e3d00000@20
  91: untyped@e3e00000@20
  92: untyped@e3f00000@20
  93: untyped@fc000000@20
  94: untyped@fc100000@20
  95: untyped@fc200000@20
  96: untyped@fc300000@20
  97: untyped@fc400000@20
  98: untyped@fc500000@20
  99: untyped@fc600000@20
  100: untyped@fc700000@20
  101: untyped@fc800000@20
  102: untyped@fc900000@20
  103: untyped@fca00000@20
  104: untyped@fcb00000@20
  105: untyped@fcc00000@20
  106: untyped@fcd00000@20
  107: untyped@fce00000@20
  108: untyped@fcf00000@20
  109: untyped@fd000000@20
  110: untyped@fd100000@20
  111: untyped@fd200000@20
  112: untyped@fd300000@20
  113: untyped@fd400000@20
  114: untyped@fd500000@20
  115: untyped@fd600000@20
  116: untyped@fd700000@20
  117: untyped@fd800000@20
  118: untyped@fd900000@20
  119: untyped@fda00000@20
  120: untyped@fdb00000@20
  121: untyped@fdc00000@20
  122: untyped@fdd00000@20
  123: untyped@fde00000@20
  124: untyped@fdf00000@20
  125: untyped@fe000000@20
  126: untyped@fe100000@20
  127: untyped@fe200000@20
  128: untyped@fe300000@20
  129: untyped@fe400000@20
  130: untyped@fe500000@20
  131: untyped@fe600000@20
  132: untyped@fe700000@20
  133: untyped@fe800000@20
  134: untyped@fe900000@20
  135: untyped@fea00000@20
  136: untyped@feb00000@20
  137: untyped@fec00000@20
  138: untyped@fed00000@20
  139: untyped@fee00000@20
  140: untyped@fef00000@20
  141: untyped@ff000000@20
  142: untyped@ff100000@20
  143: untyped@ff200000@20
  144: untyped@ff300000@20
  145: untyped@ff400000@20
  146: untyped@ff500000@20
  147: untyped@ff600000@20
  148: untyped@ff700000@20
  149: untyped@e1c00000@20
  150: untyped@e1d00000@20
  151: untyped@e1e00000@20
  152: untyped@e1f00000@20
  153: untyped@ff800000@20
  154: untyped@ff900000@20
  155: untyped@ffa00000@20
  156: untyped@ffb00000@20
  157: untyped@e0800000@20
  158: untyped@e0900000@20
  159: untyped@e0a00000@20
  160: untyped@e0b00000@20
  161: untyped@e1a00000@20
  162: untyped@e1b00000@20
  163: untyped@ffc00000@20
  164: untyped@ffd00000@20
  165: untyped@e0200000@20
  166: untyped@e0300000@20
  167: untyped@e1900000@20
  168: untyped@e8000000@20
  169: untyped@e8100000@20
  170: untyped@e8200000@20
  171: untyped@e8300000@20
  172: untyped@e8400000@20
  173: untyped@e8500000@20
  174: untyped@e8600000@20
  175: untyped@e8700000@20
  176: untyped@e8800000@20
  177: untyped@e8900000@20
  178: untyped@e8a00000@20
  179: untyped@e8b00000@20
  180: untyped@e8c00000@20
  181: untyped@e8d00000@20
  182: untyped@e8e00000@20
  183: untyped@e8f00000@20
  184: untyped@e9000000@20
  185: untyped@e9100000@20
  186: untyped@e9200000@20
  187: untyped@e9300000@20
  188: untyped@e9400000@20
  189: untyped@e9500000@20
  190: untyped@e9600000@20
  191: untyped@e9700000@20
  192: untyped@e9800000@20
  193: untyped@e9900000@20
  194: untyped@e9a00000@20
  195: untyped@e9b00000@20
  196: untyped@e9c00000@20
  197: untyped@e9d00000@20
  198: untyped@e9e00000@20
  199: untyped@e9f00000@20
  200: untyped@ea000000@20
  201: untyped@ea100000@20
  202: untyped@ea200000@20
  203: untyped@ea300000@20
  204: untyped@ea400000@20
  205: untyped@ea500000@20
  206: untyped@ea600000@20
  207: untyped@ea700000@20
  208: untyped@ea800000@20
  209: untyped@ea900000@20
  210: untyped@eaa00000@20
  211: untyped@eab00000@20
  212: untyped@eac00000@20
  213: untyped@ead00000@20
  214: untyped@eae00000@20
  215: untyped@eaf00000@20
  216: untyped@eb000000@20
  217: untyped@eb100000@20
  218: untyped@eb200000@20
  219: untyped@eb300000@20
  220: untyped@eb400000@20
  221: untyped@eb500000@20
  222: untyped@eb600000@20
  223: untyped@eb700000@20
  224: untyped@eb800000@20
  225: untyped@eb900000@20
  226: untyped@eba00000@20
  227: untyped@ebb00000@20
  228: untyped@ebc00000@20
  229: untyped@ebd00000@20
  230: untyped@ebe00000@20
  231: untyped@ebf00000@20
  232: untyped@ec000000@20
  233: untyped@ec100000@20
  234: untyped@ec200000@20
  235: untyped@ec300000@20
  236: untyped@ec400000@20
  237: untyped@ec500000@20
  238: untyped@ec600000@20
  239: untyped@ec700000@20
  240: untyped@ec800000@20
  241: untyped@ec900000@20
  242: untyped@eca00000@20
  243: untyped@ecb00000@20
  244: untyped@ecc00000@20
  245: untyped@ecd00000@20
  246: untyped@ece00000@20
  247: untyped@ecf00000@20
  248: untyped@ed000000@20
  249: untyped@ed100000@20
  250: untyped@ed200000@20
  251: untyped@ed300000@20
  252: untyped@ed400000@20
  253: untyped@ed500000@20
  254: untyped@ed600000@20
  255: untyped@ed700000@20
  256: untyped@ed800000@20
  257: untyped@ed900000@20
  258: untyped@eda00000@20
  259: untyped@edb00000@20
  260: untyped@edc00000@20
  261: untyped@edd00000@20
  262: untyped@ede00000@20
  263: untyped@edf00000@20
  264: untyped@ee000000@20
  265: untyped@ee100000@20
  266: untyped@ee200000@20
  267: untyped@ee300000@20
  268: untyped@ee400000@20
  269: untyped@ee500000@20
  270: untyped@ee600000@20
  271: untyped@ee700000@20
  272: untyped@ee800000@20
  273: untyped@ee900000@20
  274: untyped@eea00000@20
  275: untyped@eeb00000@20
  276: untyped@eec00000@20
  277: untyped@eed00000@20
  278: untyped@eee00000@20
  279: untyped@eef00000@20
  280: untyped@ef000000@20
  281: untyped@ef100000@20
  282: untyped@ef200000@20
  283: irqhandler@1b
  284: frame@d0180000
  285: frame@d0181000
  286: frame@d0182000
  287: frame@d0183000
  288: frame@d0184000
  289: frame@d0185000
  290: frame@d0186000
  291: frame@d0187000
  292: frame@d0188000
  293: frame@d0189000
  294: frame@d018a000
  295: frame@d018b000
  296: frame@d018c000
  297: frame@d018d000
  298: frame@d018e000
  299: frame@d018f000
  300: frame@d0190000
  301: frame@d0191000
  302: frame@d0192000
  303: frame@d0193000
  304: frame@d0194000
  305: frame@d0195000
  306: frame@d0196000
  307: frame@d0197000
  308: frame@d0198000
  309: frame@d0199000
  310: frame@d019a000
  311: frame@d019b000
  312: frame@d019c000
  313: frame@d019d000
  314: frame@d019e000
  315: frame@d019f000
  316: frame@d01a5000
  317: iospace@c8
  318: ep@e001cff0 ( W )
  319: aep@fffeffd0 (badge: 0x0,  R)
}
cnode@f6bcc000{
  0: cnode@f6bc8000
}
pd@f6c7f000{
  0x0: pt@f6dff000
  0x340: pt@f6df5000
}
pd@f6c7e000{
  0x0: pt@f6dfd000
  0x300: pt@f6df9000
  0x340: pt@f6df4000
}
pd@f6c7d000{
  0x0: pt@f6dfc000
  0x1: pt@f6dfb000
  0x340: pt@f6dfa000
}
pd@f6c7c000{
  0x0: pt@f6df8000
  0x1: pt@f6df7000
  0x300: pt@f6df6000
  0x340: pt@f6df3000
}
pt@f6df5000{
  0x0: frame@f6cff000(RW)
  0x1: frame@f9dc7000(RW)
  0x2: frame@f9dc8000(RW)
}
pt@f6dff000{
  0x10: frame@f6cfe000(R )
  0x11: frame@f6cfd000(R )
  0x12: frame@f6cfc000(R )
  0x13: frame@f6cfb000(R )
  0x14: frame@f6cfa000(R )
  0x15: frame@f6cf9000(RW)
  0x16: frame@f6cf8000(RW)
  0x17: frame@f6cf7000(RW)
  0x18: frame@f6cf6000(RW)
  0x19: frame@f6cf5000(RW)
  0x1a: frame@f6cf4000(RW)
  0x1b: frame@f6cf3000(RW)
  0x1c: frame@f6cf2000(RW)
}
pt@f6df4000{
  0x0: frame@f6cf1000(RW)
  0x1: frame@f9dc5000(RW)
  0x2: frame@f9dc6000(RW)
}
pt@f6df9000{
  0x200: frame@d0200000(RW)
  0x201: frame@d0201000(RW)
  0x202: frame@d0202000(RW)
  0x203: frame@d0203000(RW)
  0x204: frame@d0204000(RW)
  0x205: frame@d0205000(RW)
  0x206: frame@d0206000(RW)
  0x207: frame@d0207000(RW)
  0x208: frame@d0208000(RW)
  0x209: frame@d0209000(RW)
  0x20a: frame@d020a000(RW)
  0x20b: frame@d020b000(RW)
  0x20c: frame@d020c000(RW)
  0x20d: frame@d020d000(RW)
  0x20e: frame@d020e000(RW)
  0x20f: frame@d020f000(RW)
  0x210: frame@d0210000(RW)
  0x211: frame@d0211000(RW)
  0x212: frame@d0212000(RW)
  0x213: frame@d0213000(RW)
  0x214: frame@d0214000(RW)
  0x215: frame@d0215000(RW)
  0x216: frame@d0216000(RW)
  0x217: frame@d0217000(RW)
  0x218: frame@d0218000(RW)
  0x219: frame@d0219000(RW)
  0x21a: frame@d021a000(RW)
  0x21b: frame@d021b000(RW)
  0x21c: frame@d021c000(RW)
  0x21d: frame@d021d000(RW)
  0x21e: frame@d021e000(RW)
  0x21f: frame@d021f000(RW)
  0x220: frame@d0220000(RW)
  0x221: frame@d0221000(RW)
  0x222: frame@d0222000(RW)
  0x223: frame@d0223000(RW)
  0x224: frame@d0224000(RW)
  0x225: frame@d0225000(RW)
  0x226: frame@d0226000(RW)
  0x227: frame@d0227000(RW)
  0x228: frame@d0228000(RW)
  0x229: frame@d0229000(RW)
  0x22a: frame@d022a000(RW)
  0x22b: frame@d022b000(RW)
  0x22c: frame@d022c000(RW)
  0x22d: frame@d022d000(RW)
  0x22e: frame@d022e000(RW)
  0x22f: frame@d022f000(RW)
  0x230: frame@d0230000(RW)
  0x231: frame@d0231000(RW)
  0x232: frame@d0232000(RW)
  0x233: frame@d0233000(RW)
  0x234: frame@d0234000(RW)
  0x235: frame@d0235000(RW)
  0x236: frame@d0236000(RW)
  0x237: frame@d0237000(RW)
  0x238: frame@d0238000(RW)
  0x239: frame@d0239000(RW)
  0x23a: frame@d023a000(RW)
  0x23b: frame@d023b000(RW)
  0x23c: frame@d023c000(RW)
  0x23d: frame@d023d000(RW)
  0x23e: frame@d023e000(RW)
  0x23f: frame@d023f000(RW)
  0x240: frame@d0240000(RW)
  0x241: frame@d0241000(RW)
  0x242: frame@d0242000(RW)
  0x243: frame@d0243000(RW)
  0x244: frame@d0244000(RW)
  0x245: frame@d0245000(RW)
  0x246: frame@d0246000(RW)
  0x247: frame@d0247000(RW)
  0x248: frame@d0248000(RW)
  0x249: frame@d0249000(RW)
  0x24a: frame@d024a000(RW)
  0x24b: frame@d024b000(RW)
  0x24c: frame@d024c000(RW)
  0x24d: frame@d024d000(RW)
  0x24e: frame@d024e000(RW)
  0x24f: frame@d024f000(RW)
  0x250: frame@d0250000(RW)
  0x251: frame@d0251000(RW)
  0x252: frame@d0252000(RW)
  0x253: frame@d0253000(RW)
  0x254: frame@d0254000(RW)
  0x255: frame@d0255000(RW)
  0x256: frame@d0256000(RW)
  0x257: frame@d0257000(RW)
  0x258: frame@d0258000(RW)
  0x259: frame@d0259000(RW)
  0x25a: frame@d025a000(RW)
  0x25b: frame@d025b000(RW)
  0x25c: frame@d025c000(RW)
  0x25d: frame@d025d000(RW)
  0x25e: frame@d025e000(RW)
  0x25f: frame@d025f000(RW)
  0x260: frame@d0260000(RW)
  0x261: frame@d0261000(RW)
  0x262: frame@d0262000(RW)
  0x263: frame@d0263000(RW)
  0x264: frame@d0264000(RW)
  0x265: frame@d0265000(RW)
  0x266: frame@d0266000(RW)
  0x267: frame@d0267000(RW)
  0x268: frame@d0268000(RW)
  0x269: frame@d0269000(RW)
  0x26a: frame@d026a000(RW)
  0x26b: frame@d026b000(RW)
  0x26c: frame@d026c000(RW)
  0x26d: frame@d026d000(RW)
  0x26e: frame@d026e000(RW)
  0x26f: frame@d026f000(RW)
  0x270: frame@d0270000(RW)
  0x271: frame@d0271000(RW)
  0x272: frame@d0272000(RW)
  0x273: frame@d0273000(RW)
  0x274: frame@d0274000(RW)
  0x275: frame@d0275000(RW)
  0x276: frame@d0276000(RW)
  0x277: frame@d0277000(RW)
  0x278: frame@d0278000(RW)
  0x279: frame@d0279000(RW)
  0x27a: frame@d027a000(RW)
  0x27b: frame@d027b000(RW)
  0x27c: frame@d027c000(RW)
  0x27d: frame@d027d000(RW)
  0x27e: frame@d027e000(RW)
  0x27f: frame@d027f000(RW)
  0x300: frame@d0300000(RW)
  0x301: frame@d0301000(RW)
  0x302: frame@d0302000(RW)
  0x303: frame@d0303000(RW)
}
pt@f6dfd000{
  0x10: frame@f6cf0000(R )
  0x11: frame@f6cef000(R )
  0x12: frame@f6cee000(R )
  0x13: frame@f6ced000(R )
  0x14: frame@f6cec000(RW)
  0x15: frame@f6ceb000(RW)
  0x16: frame@f6cea000(RW)
}
pt@f6dfa000{
  0x0: frame@f729e000(R )
  0x1: frame@f9dc4000(R )
}
pt@f6dfb000{
  0x0: frame@f71f9000(R )
  0x1: frame@f71f8000(R )
  0x2: frame@f71f7000(R )
  0x3: frame@f71f6000(R )
  0x4: frame@f71f5000(R )
  0x5: frame@f71f4000(R )
  0x6: frame@f71f3000(R )
  0x7: frame@f71f2000(R )
  0x8: frame@f71f1000(R )
  0x9: frame@f71f0000(R )
  0xa: frame@f71ef000(R )
  0xb: frame@f71ee000(R )
  0xc: frame@f71ed000(R )
  0xd: frame@f71ec000(R )
  0xe: frame@f71eb000(R )
  0xf: frame@f71ea000(R )
  0x10: frame@f71e9000(R )
  0x11: frame@f71e8000(R )
  0x12: frame@f71e7000(R )
  0x13: frame@f71e6000(R )
  0x14: frame@f71e5000(R )
  0x15: frame@f71e4000(R )
  0x16: frame@f71e3000(R )
  0x17: frame@f71e2000(R )
  0x18: frame@f71e1000(R )
  0x19: frame@f71e0000(R )
  0x1a: frame@f71df000(R )
  0x1b: frame@f71de000(R )
  0x1c: frame@f71dd000(R )
  0x1d: frame@f71dc000(R )
  0x1e: frame@f71db000(R )
  0x1f: frame@f71da000(R )
  0x20: frame@f71d9000(R )
  0x21: frame@f71d8000(R )
  0x22: frame@f71d7000(R )
  0x23: frame@f71d6000(R )
  0x24: frame@f71d5000(R )
  0x25: frame@f71d4000(R )
  0x26: frame@f71d3000(R )
  0x27: frame@f71d2000(R )
  0x28: frame@f71d1000(R )
  0x29: frame@f71d0000(R )
  0x2a: frame@f71cf000(R )
  0x2b: frame@f71ce000(R )
  0x2c: frame@f71cd000(R )
  0x2d: frame@f71cc000(R )
  0x2e: frame@f71cb000(R )
  0x2f: frame@f71ca000(R )
  0x30: frame@f71c9000(R )
  0x31: frame@f71c8000(R )
  0x32: frame@f71c7000(R )
  0x33: frame@f71c6000(R )
  0x34: frame@f71c5000(R )
  0x35: frame@f71c4000(R )
  0x36: frame@f71c3000(R )
  0x37: frame@f71c2000(R )
  0x38: frame@f71c1000(R )
  0x39: frame@f71c0000(R )
  0x3a: frame@f71bf000(R )
  0x3b: frame@f71be000(R )
  0x3c: frame@f71bd000(R )
  0x3d: frame@f71bc000(R )
  0x3e: frame@f71bb000(R )
  0x3f: frame@f71ba000(R )
  0x40: frame@f71b9000(R )
  0x41: frame@f71b8000(R )
  0x42: frame@f71b7000(R )
  0x43: frame@f71b6000(R )
  0x44: frame@f71b5000(R )
  0x45: frame@f71b4000(R )
  0x46: frame@f71b3000(R )
  0x47: frame@f71b2000(R )
  0x48: frame@f71b1000(R )
  0x49: frame@f71b0000(R )
  0x4a: frame@f71af000(R )
  0x4b: frame@f71ae000(R )
  0x4c: frame@f71ad000(R )
  0x4d: frame@f71ac000(R )
  0x4e: frame@f71ab000(R )
  0x4f: frame@f71aa000(R )
  0x50: frame@f71a9000(R )
  0x51: frame@f71a8000(R )
  0x52: frame@f71a7000(R )
  0x53: frame@f71a6000(R )
  0x54: frame@f71a5000(R )
  0x55: frame@f71a4000(R )
  0x56: frame@f71a3000(R )
  0x57: frame@f71a2000(R )
  0x58: frame@f71a1000(R )
  0x59: frame@f71a0000(R )
  0x5a: frame@f719f000(R )
  0x5b: frame@f719e000(R )
  0x5c: frame@f719d000(R )
  0x5d: frame@f719c000(R )
  0x5e: frame@f719b000(R )
  0x5f: frame@f719a000(R )
  0x60: frame@f7199000(R )
  0x61: frame@f7198000(R )
  0x62: frame@f7197000(R )
  0x63: frame@f7196000(R )
  0x64: frame@f7195000(R )
  0x65: frame@f7194000(R )
  0x66: frame@f7193000(R )
  0x67: frame@f7192000(R )
  0x68: frame@f7191000(R )
  0x69: frame@f7190000(R )
  0x6a: frame@f718f000(R )
  0x6b: frame@f718e000(R )
  0x6c: frame@f718d000(R )
  0x6d: frame@f718c000(R )
  0x6e: frame@f718b000(R )
  0x6f: frame@f718a000(R )
  0x70: frame@f7189000(R )
  0x71: frame@f7188000(R )
  0x72: frame@f7187000(R )
  0x73: frame@f7186000(R )
  0x74: frame@f7185000(R )
  0x75: frame@f7184000(R )
  0x76: frame@f7183000(R )
  0x77: frame@f7182000(R )
  0x78: frame@f7181000(R )
  0x79: frame@f7180000(R )
  0x7a: frame@f717f000(R )
  0x7b: frame@f717e000(R )
  0x7c: frame@f717d000(R )
  0x7d: frame@f717c000(R )
  0x7e: frame@f717b000(R )
  0x7f: frame@f717a000(R )
  0x80: frame@f7179000(R )
  0x81: frame@f7178000(R )
  0x82: frame@f7177000(R )
  0x83: frame@f7176000(R )
  0x84: frame@f7175000(R )
  0x85: frame@f7174000(R )
  0x86: frame@f7173000(R )
  0x87: frame@f7172000(R )
  0x88: frame@f7171000(R )
  0x89: frame@f7170000(R )
  0x8a: frame@f716f000(R )
  0x8b: frame@f716e000(R )
  0x8c: frame@f716d000(R )
  0x8d: frame@f716c000(R )
  0x8e: frame@f716b000(R )
  0x8f: frame@f716a000(R )
  0x90: frame@f7169000(R )
  0x91: frame@f7168000(R )
  0x92: frame@f7167000(R )
  0x93: frame@f7166000(R )
  0x94: frame@f7165000(R )
  0x95: frame@f7164000(R )
  0x96: frame@f7163000(R )
  0x97: frame@f7162000(R )
  0x98: frame@f7161000(R )
  0x99: frame@f7160000(R )
  0x9a: frame@f715f000(R )
  0x9b: frame@f715e000(R )
  0x9c: frame@f715d000(R )
  0x9d: frame@f715c000(R )
  0x9e: frame@f715b000(R )
  0x9f: frame@f715a000(R )
  0xa0: frame@f7159000(R )
  0xa1: frame@f7158000(R )
  0xa2: frame@f7157000(R )
  0xa3: frame@f7156000(R )
  0xa4: frame@f7155000(R )
  0xa5: frame@f7154000(R )
  0xa6: frame@f7153000(R )
  0xa7: frame@f7152000(R )
  0xa8: frame@f7151000(R )
  0xa9: frame@f7150000(R )
  0xaa: frame@f714f000(R )
  0xab: frame@f714e000(R )
  0xac: frame@f714d000(R )
  0xad: frame@f714c000(R )
  0xae: frame@f714b000(R )
  0xaf: frame@f714a000(R )
  0xb0: frame@f7149000(R )
  0xb1: frame@f7148000(R )
  0xb2: frame@f7147000(R )
  0xb3: frame@f7146000(R )
  0xb4: frame@f7145000(R )
  0xb5: frame@f7144000(R )
  0xb6: frame@f7143000(R )
  0xb7: frame@f7142000(R )
  0xb8: frame@f7141000(R )
  0xb9: frame@f7140000(R )
  0xba: frame@f713f000(R )
  0xbb: frame@f713e000(R )
  0xbc: frame@f713d000(R )
  0xbd: frame@f713c000(R )
  0xbe: frame@f713b000(R )
  0xbf: frame@f713a000(R )
  0xc0: frame@f7139000(R )
  0xc1: frame@f7138000(R )
  0xc2: frame@f7137000(R )
  0xc3: frame@f7136000(R )
  0xc4: frame@f7135000(R )
  0xc5: frame@f7134000(R )
  0xc6: frame@f7133000(R )
  0xc7: frame@f7132000(R )
  0xc8: frame@f7131000(R )
  0xc9: frame@f7130000(R )
  0xca: frame@f712f000(R )
  0xcb: frame@f712e000(R )
  0xcc: frame@f712d000(R )
  0xcd: frame@f712c000(R )
  0xce: frame@f712b000(R )
  0xcf: frame@f712a000(R )
  0xd0: frame@f7129000(R )
  0xd1: frame@f7128000(R )
  0xd2: frame@f7127000(R )
  0xd3: frame@f7126000(R )
  0xd4: frame@f7125000(R )
  0xd5: frame@f7124000(R )
  0xd6: frame@f7123000(R )
  0xd7: frame@f7122000(R )
  0xd8: frame@f7121000(R )
  0xd9: frame@f7120000(R )
  0xda: frame@f711f000(R )
  0xdb: frame@f711e000(R )
  0xdc: frame@f711d000(R )
  0xdd: frame@f711c000(R )
  0xde: frame@f711b000(R )
  0xdf: frame@f711a000(R )
  0xe0: frame@f7119000(R )
  0xe1: frame@f7118000(R )
  0xe2: frame@f7117000(R )
  0xe3: frame@f7116000(R )
  0xe4: frame@f7115000(R )
  0xe5: frame@f7114000(R )
  0xe6: frame@f7113000(R )
  0xe7: frame@f7112000(R )
  0xe8: frame@f7111000(R )
  0xe9: frame@f7110000(R )
  0xea: frame@f710f000(R )
  0xeb: frame@f710e000(R )
  0xec: frame@f710d000(R )
  0xed: frame@f710c000(R )
  0xee: frame@f710b000(R )
  0xef: frame@f710a000(R )
  0xf0: frame@f7109000(R )
  0xf1: frame@f7108000(R )
  0xf2: frame@f7107000(R )
  0xf3: frame@f7106000(R )
  0xf4: frame@f7105000(R )
  0xf5: frame@f7104000(R )
  0xf6: frame@f7103000(R )
  0xf7: frame@f7102000(R )
  0xf8: frame@f7101000(R )
  0xf9: frame@f7100000(R )
  0xfa: frame@f72ff000(R )
  0xfb: frame@f72fe000(R )
  0xfc: frame@f72fd000(R )
  0xfd: frame@f72fc000(R )
  0xfe: frame@f72fb000(R )
  0xff: frame@f72fa000(R )
  0x100: frame@f72f9000(R )
  0x101: frame@f72f8000(R )
  0x102: frame@f72f7000(R )
  0x103: frame@f72f6000(R )
  0x104: frame@f72f5000(R )
  0x105: frame@f72f4000(R )
  0x106: frame@f72f3000(R )
  0x107: frame@f72f2000(R )
  0x108: frame@f72f1000(R )
  0x109: frame@f72f0000(R )
  0x10a: frame@f72ef000(R )
  0x10b: frame@f72ee000(R )
  0x10c: frame@f72ed000(R )
  0x10d: frame@f72ec000(R )
  0x10e: frame@f72eb000(R )
  0x10f: frame@f72ea000(R )
  0x110: frame@f72e9000(R )
  0x111: frame@f72e8000(R )
  0x112: frame@f72e7000(R )
  0x113: frame@f72e6000(R )
  0x114: frame@f72e5000(R )
  0x115: frame@f72e4000(R )
  0x116: frame@f72e3000(R )
  0x117: frame@f72e2000(R )
  0x118: frame@f72e1000(R )
  0x119: frame@f72e0000(R )
  0x11a: frame@f72df000(R )
  0x11b: frame@f72de000(R )
  0x11c: frame@f72dd000(R )
  0x11d: frame@f72dc000(R )
  0x11e: frame@f72db000(R )
  0x11f: frame@f72da000(R )
  0x120: frame@f72d9000(R )
  0x121: frame@f72d8000(R )
  0x122: frame@f72d7000(R )
  0x123: frame@f72d6000(R )
  0x124: frame@f72d5000(R )
  0x125: frame@f72d4000(R )
  0x126: frame@f72d3000(R )
  0x127: frame@f72d2000(R )
  0x128: frame@f72d1000(R )
  0x129: frame@f72d0000(R )
  0x12a: frame@f72cf000(R )
  0x12b: frame@f72ce000(R )
  0x12c: frame@f72cd000(R )
  0x12d: frame@f72cc000(R )
  0x12e: frame@f72cb000(R )
  0x12f: frame@f72ca000(R )
  0x130: frame@f72c9000(R )
  0x131: frame@f72c8000(R )
  0x132: frame@f72c7000(R )
  0x133: frame@f72c6000(R )
  0x134: frame@f72c5000(R )
  0x135: frame@f72c4000(R )
  0x136: frame@f72c3000(R )
  0x137: frame@f72c2000(R )
  0x138: frame@f72c1000(R )
  0x139: frame@f72c0000(R )
  0x13a: frame@f72bf000(R )
  0x13b: frame@f72be000(R )
  0x13c: frame@f72bd000(R )
  0x13d: frame@f72bc000(R )
  0x13e: frame@f72bb000(R )
  0x13f: frame@f72ba000(R )
  0x140: frame@f72b9000(R )
  0x141: frame@f72b8000(R )
  0x142: frame@f72b7000(R )
  0x143: frame@f72b6000(R )
  0x144: frame@f72b5000(R )
  0x145: frame@f72b4000(R )
  0x146: frame@f72b3000(R )
  0x147: frame@f72b2000(R )
  0x148: frame@f72b1000(R )
  0x149: frame@f72b0000(R )
  0x14a: frame@f72af000(R )
  0x14b: frame@f72ae000(R )
  0x14c: frame@f72ad000(R )
  0x14d: frame@f72ac000(R )
  0x14e: frame@f72ab000(R )
  0x14f: frame@f72aa000(R )
  0x150: frame@f72a9000(R )
  0x151: frame@f72a8000(R )
  0x152: frame@f72a7000(R )
  0x153: frame@f72a6000(R )
  0x154: frame@f72a5000(R )
  0x155: frame@f72a4000(R )
  0x156: frame@f72a3000(R )
  0x157: frame@f72a2000(R )
  0x158: frame@f72a1000(R )
  0x159: frame@f72a0000(R )
  0x15a: frame@f729f000(R )
}
pt@f6dfc000{
  0x10: frame@f6ce9000(R )
  0x11: frame@f6ce8000(R )
  0x12: frame@f6ce7000(R )
  0x13: frame@f6ce6000(R )
  0x14: frame@f6ce5000(R )
  0x15: frame@f6ce4000(R )
  0x16: frame@f6ce3000(R )
  0x17: frame@f6ce2000(R )
  0x18: frame@f6ce1000(R )
  0x19: frame@f6ce0000(R )
  0x1a: frame@f6cdf000(R )
  0x1b: frame@f6cde000(R )
  0x1c: frame@f6cdd000(R )
  0x1d: frame@f6cdc000(R )
  0x1e: frame@f6cdb000(R )
  0x1f: frame@f6cda000(R )
  0x20: frame@f6cd9000(R )
  0x21: frame@f6cd8000(R )
  0x22: frame@f6cd7000(R )
  0x23: frame@f6cd6000(R )
  0x24: frame@f6cd5000(R )
  0x25: frame@f6cd4000(R )
  0x26: frame@f6cd3000(R )
  0x27: frame@f6cd2000(R )
  0x28: frame@f6cd1000(R )
  0x29: frame@f6cd0000(R )
  0x2a: frame@f6ccf000(R )
  0x2b: frame@f6cce000(R )
  0x2c: frame@f6ccd000(R )
  0x2d: frame@f6ccc000(R )
  0x2e: frame@f6ccb000(R )
  0x2f: frame@f6cca000(R )
  0x30: frame@f6cc9000(R )
  0x31: frame@f6cc8000(R )
  0x32: frame@f6cc7000(R )
  0x33: frame@f6cc6000(R )
  0x34: frame@f6cc5000(R )
  0x35: frame@f6cc4000(R )
  0x36: frame@f6cc3000(R )
  0x37: frame@f6cc2000(R )
  0x38: frame@f6cc1000(R )
  0x39: frame@f6cc0000(R )
  0x3a: frame@f6cbf000(R )
  0x3b: frame@f6cbe000(R )
  0x3c: frame@f6cbd000(R )
  0x3d: frame@f6cbc000(R )
  0x3e: frame@f6cbb000(R )
  0x3f: frame@f6cba000(R )
  0x40: frame@f6cb9000(R )
  0x41: frame@f6cb8000(R )
  0x42: frame@f6cb7000(R )
  0x43: frame@f6cb6000(R )
  0x44: frame@f6cb5000(R )
  0x45: frame@f6cb4000(R )
  0x46: frame@f6cb3000(R )
  0x47: frame@f6cb2000(R )
  0x48: frame@f6cb1000(R )
  0x49: frame@f6cb0000(R )
  0x4a: frame@f6caf000(R )
  0x4b: frame@f6cae000(R )
  0x4c: frame@f6cad000(R )
  0x4d: frame@f6cac000(R )
  0x4e: frame@f6cab000(R )
  0x4f: frame@f6caa000(R )
  0x50: frame@f6ca9000(R )
  0x51: frame@f6ca8000(R )
  0x52: frame@f6ca7000(R )
  0x53: frame@f6ca6000(R )
  0x54: frame@f6ca5000(R )
  0x55: frame@f6ca4000(R )
  0x56: frame@f6ca3000(R )
  0x57: frame@f6ca2000(R )
  0x58: frame@f6ca1000(R )
  0x59: frame@f6ca0000(R )
  0x5a: frame@f6c9f000(R )
  0x5b: frame@f6c9e000(R )
  0x5c: frame@f6c9d000(R )
  0x5d: frame@f6c9c000(R )
  0x5e: frame@f6c9b000(R )
  0x5f: frame@f6c9a000(R )
  0x60: frame@f6c99000(R )
  0x61: frame@f6c98000(R )
  0x62: frame@f6c97000(R )
  0x63: frame@f6c96000(R )
  0x64: frame@f6c95000(R )
  0x65: frame@f6c94000(R )
  0x66: frame@f6c93000(R )
  0x67: frame@f6c92000(R )
  0x68: frame@f6c91000(R )
  0x69: frame@f6c90000(R )
  0x6a: frame@f6c8f000(R )
  0x6b: frame@f6c8e000(R )
  0x6c: frame@f6c8d000(R )
  0x6d: frame@f6c8c000(R )
  0x6e: frame@f6c8b000(R )
  0x6f: frame@f6c8a000(R )
  0x70: frame@f6c89000(R )
  0x71: frame@f6c88000(R )
  0x72: frame@f6c87000(R )
  0x73: frame@f6c86000(R )
  0x74: frame@f6c85000(R )
  0x75: frame@f6c84000(R )
  0x76: frame@f6c83000(R )
  0x77: frame@f6c82000(R )
  0x78: frame@f6c81000(R )
  0x79: frame@f6c80000(R )
  0x7a: frame@f6d7f000(R )
  0x7b: frame@f6d7e000(R )
  0x7c: frame@f6d7d000(R )
  0x7d: frame@f6d7c000(R )
  0x7e: frame@f6d7b000(R )
  0x7f: frame@f6d7a000(R )
  0x80: frame@f6d79000(R )
  0x81: frame@f6d78000(R )
  0x82: frame@f6d77000(R )
  0x83: frame@f6d76000(R )
  0x84: frame@f6d75000(R )
  0x85: frame@f6d74000(R )
  0x86: frame@f6d73000(R )
  0x87: frame@f6d72000(R )
  0x88: frame@f6d71000(R )
  0x89: frame@f6d70000(R )
  0x8a: frame@f6d6f000(R )
  0x8b: frame@f6d6e000(R )
  0x8c: frame@f6d6d000(R )
  0x8d: frame@f6d6c000(R )
  0x8e: frame@f6d6b000(R )
  0x8f: frame@f6d6a000(R )
  0x90: frame@f6d69000(R )
  0x91: frame@f6d68000(R )
  0x92: frame@f6d67000(R )
  0x93: frame@f6d66000(R )
  0x94: frame@f6d65000(R )
  0x95: frame@f6d64000(R )
  0x96: frame@f6d63000(R )
  0x97: frame@f6d62000(R )
  0x98: frame@f6d61000(R )
  0x99: frame@f6d60000(R )
  0x9a: frame@f6d5f000(R )
  0x9b: frame@f6d5e000(R )
  0x9c: frame@f6d5d000(R )
  0x9d: frame@f6d5c000(R )
  0x9e: frame@f6d5b000(R )
  0x9f: frame@f6d5a000(R )
  0xa0: frame@f6d59000(R )
  0xa1: frame@f6d58000(R )
  0xa2: frame@f6d57000(R )
  0xa3: frame@f6d56000(R )
  0xa4: frame@f6d55000(R )
  0xa5: frame@f6d54000(R )
  0xa6: frame@f6d53000(R )
  0xa7: frame@f6d52000(R )
  0xa8: frame@f6d51000(R )
  0xa9: frame@f6d50000(R )
  0xaa: frame@f6d4f000(R )
  0xab: frame@f6d4e000(R )
  0xac: frame@f6d4d000(R )
  0xad: frame@f6d4c000(R )
  0xae: frame@f6d4b000(R )
  0xaf: frame@f6d4a000(R )
  0xb0: frame@f6d49000(R )
  0xb1: frame@f6d48000(R )
  0xb2: frame@f6d47000(R )
  0xb3: frame@f6d46000(R )
  0xb4: frame@f6d45000(R )
  0xb5: frame@f6d44000(R )
  0xb6: frame@f6d43000(R )
  0xb7: frame@f6d42000(R )
  0xb8: frame@f6d41000(R )
  0xb9: frame@f6d40000(R )
  0xba: frame@f6d3f000(R )
  0xbb: frame@f6d3e000(R )
  0xbc: frame@f6d3d000(R )
  0xbd: frame@f6d3c000(R )
  0xbe: frame@f6d3b000(R )
  0xbf: frame@f6d3a000(R )
  0xc0: frame@f6d39000(R )
  0xc1: frame@f6d38000(R )
  0xc2: frame@f6d37000(R )
  0xc3: frame@f6d36000(R )
  0xc4: frame@f6d35000(R )
  0xc5: frame@f6d34000(R )
  0xc6: frame@f6d33000(R )
  0xc7: frame@f6d32000(R )
  0xc8: frame@f6d31000(R )
  0xc9: frame@f6d30000(R )
  0xca: frame@f6d2f000(R )
  0xcb: frame@f6d2e000(R )
  0xcc: frame@f6d2d000(R )
  0xcd: frame@f6d2c000(R )
  0xce: frame@f6d2b000(R )
  0xcf: frame@f6d2a000(R )
  0xd0: frame@f6d29000(R )
  0xd1: frame@f6d28000(R )
  0xd2: frame@f6d27000(R )
  0xd3: frame@f6d26000(R )
  0xd4: frame@f6d25000(R )
  0xd5: frame@f6d24000(R )
  0xd6: frame@f6d23000(R )
  0xd7: frame@f6d22000(R )
  0xd8: frame@f6d21000(R )
  0xd9: frame@f6d20000(R )
  0xda: frame@f6d1f000(R )
  0xdb: frame@f6d1e000(R )
  0xdc: frame@f6d1d000(R )
  0xdd: frame@f6d1c000(R )
  0xde: frame@f6d1b000(R )
  0xdf: frame@f6d1a000(R )
  0xe0: frame@f6d19000(R )
  0xe1: frame@f6d18000(R )
  0xe2: frame@f6d17000(R )
  0xe3: frame@f6d16000(R )
  0xe4: frame@f6d15000(R )
  0xe5: frame@f6d14000(R )
  0xe6: frame@f6d13000(R )
  0xe7: frame@f6d12000(R )
  0xe8: frame@f6d11000(R )
  0xe9: frame@f6d10000(R )
  0xea: frame@f6d0f000(R )
  0xeb: frame@f6d0e000(R )
  0xec: frame@f6d0d000(R )
  0xed: frame@f6d0c000(R )
  0xee: frame@f6d0b000(R )
  0xef: frame@f6d0a000(R )
  0xf0: frame@f6d09000(R )
  0xf1: frame@f6d08000(R )
  0xf2: frame@f6d07000(R )
  0xf3: frame@f6d06000(R )
  0xf4: frame@f6d05000(R )
  0xf5: frame@f6d04000(R )
  0xf6: frame@f6d03000(R )
  0xf7: frame@f6d02000(R )
  0xf8: frame@f6d01000(R )
  0xf9: frame@f6d00000(R )
  0xfa: frame@f6eff000(R )
  0xfb: frame@f6efe000(R )
  0xfc: frame@f6efd000(R )
  0xfd: frame@f6efc000(R )
  0xfe: frame@f6efb000(R )
  0xff: frame@f6efa000(R )
  0x100: frame@f6ef9000(R )
  0x101: frame@f6ef8000(R )
  0x102: frame@f6ef7000(R )
  0x103: frame@f6ef6000(R )
  0x104: frame@f6ef5000(R )
  0x105: frame@f6ef4000(R )
  0x106: frame@f6ef3000(R )
  0x107: frame@f6ef2000(R )
  0x108: frame@f6ef1000(R )
  0x109: frame@f6ef0000(R )
  0x10a: frame@f6eef000(R )
  0x10b: frame@f6eee000(R )
  0x10c: frame@f6eed000(R )
  0x10d: frame@f6eec000(R )
  0x10e: frame@f6eeb000(R )
  0x10f: frame@f6eea000(R )
  0x110: frame@f6ee9000(R )
  0x111: frame@f6ee8000(R )
  0x112: frame@f6ee7000(R )
  0x113: frame@f6ee6000(R )
  0x114: frame@f6ee5000(R )
  0x115: frame@f6ee4000(R )
  0x116: frame@f6ee3000(R )
  0x117: frame@f6ee2000(R )
  0x118: frame@f6ee1000(R )
  0x119: frame@f6ee0000(R )
  0x11a: frame@f6edf000(R )
  0x11b: frame@f6ede000(R )
  0x11c: frame@f6edd000(R )
  0x11d: frame@f6edc000(R )
  0x11e: frame@f6edb000(R )
  0x11f: frame@f6eda000(R )
  0x120: frame@f6ed9000(R )
  0x121: frame@f6ed8000(R )
  0x122: frame@f6ed7000(R )
  0x123: frame@f6ed6000(R )
  0x124: frame@f6ed5000(R )
  0x125: frame@f6ed4000(R )
  0x126: frame@f6ed3000(R )
  0x127: frame@f6ed2000(R )
  0x128: frame@f6ed1000(R )
  0x129: frame@f6ed0000(R )
  0x12a: frame@f6ecf000(R )
  0x12b: frame@f6ece000(R )
  0x12c: frame@f6ecd000(R )
  0x12d: frame@f6ecc000(R )
  0x12e: frame@f6ecb000(R )
  0x12f: frame@f6eca000(R )
  0x130: frame@f6ec9000(R )
  0x131: frame@f6ec8000(R )
  0x132: frame@f6ec7000(R )
  0x133: frame@f6ec6000(R )
  0x134: frame@f6ec5000(R )
  0x135: frame@f6ec4000(R )
  0x136: frame@f6ec3000(R )
  0x137: frame@f6ec2000(R )
  0x138: frame@f6ec1000(R )
  0x139: frame@f6ec0000(R )
  0x13a: frame@f6ebf000(R )
  0x13b: frame@f6ebe000(R )
  0x13c: frame@f6ebd000(R )
  0x13d: frame@f6ebc000(R )
  0x13e: frame@f6ebb000(R )
  0x13f: frame@f6eba000(R )
  0x140: frame@f6eb9000(R )
  0x141: frame@f6eb8000(R )
  0x142: frame@f6eb7000(R )
  0x143: frame@f6eb6000(R )
  0x144: frame@f6eb5000(R )
  0x145: frame@f6eb4000(R )
  0x146: frame@f6eb3000(R )
  0x147: frame@f6eb2000(R )
  0x148: frame@f6eb1000(R )
  0x149: frame@f6eb0000(R )
  0x14a: frame@f6eaf000(R )
  0x14b: frame@f6eae000(R )
  0x14c: frame@f6ead000(R )
  0x14d: frame@f6eac000(R )
  0x14e: frame@f6eab000(R )
  0x14f: frame@f6eaa000(R )
  0x150: frame@f6ea9000(R )
  0x151: frame@f6ea8000(R )
  0x152: frame@f6ea7000(R )
  0x153: frame@f6ea6000(R )
  0x154: frame@f6ea5000(R )
  0x155: frame@f6ea4000(R )
  0x156: frame@f6ea3000(R )
  0x157: frame@f6ea2000(R )
  0x158: frame@f6ea1000(R )
  0x159: frame@f6ea0000(R )
  0x15a: frame@f6e9f000(R )
  0x15b: frame@f6e9e000(R )
  0x15c: frame@f6e9d000(R )
  0x15d: frame@f6e9c000(R )
  0x15e: frame@f6e9b000(R )
  0x15f: frame@f6e9a000(R )
  0x160: frame@f6e99000(R )
  0x161: frame@f6e98000(R )
  0x162: frame@f6e97000(R )
  0x163: frame@f6e96000(R )
  0x164: frame@f6e95000(R )
  0x165: frame@f6e94000(R )
  0x166: frame@f6e93000(R )
  0x167: frame@f6e92000(R )
  0x168: frame@f6e91000(R )
  0x169: frame@f6e90000(R )
  0x16a: frame@f6e8f000(R )
  0x16b: frame@f6e8e000(R )
  0x16c: frame@f6e8d000(R )
  0x16d: frame@f6e8c000(R )
  0x16e: frame@f6e8b000(R )
  0x16f: frame@f6e8a000(R )
  0x170: frame@f6e89000(R )
  0x171: frame@f6e88000(R )
  0x172: frame@f6e87000(R )
  0x173: frame@f6e86000(R )
  0x174: frame@f6e85000(R )
  0x175: frame@f6e84000(R )
  0x176: frame@f6e83000(R )
  0x177: frame@f6e82000(R )
  0x178: frame@f6e81000(R )
  0x179: frame@f6e80000(R )
  0x17a: frame@f6e7f000(R )
  0x17b: frame@f6e7e000(R )
  0x17c: frame@f6e7d000(R )
  0x17d: frame@f6e7c000(R )
  0x17e: frame@f6e7b000(R )
  0x17f: frame@f6e7a000(R )
  0x180: frame@f6e79000(R )
  0x181: frame@f6e78000(R )
  0x182: frame@f6e77000(R )
  0x183: frame@f6e76000(R )
  0x184: frame@f6e75000(R )
  0x185: frame@f6e74000(R )
  0x186: frame@f6e73000(R )
  0x187: frame@f6e72000(R )
  0x188: frame@f6e71000(R )
  0x189: frame@f6e70000(R )
  0x18a: frame@f6e6f000(R )
  0x18b: frame@f6e6e000(R )
  0x18c: frame@f6e6d000(R )
  0x18d: frame@f6e6c000(R )
  0x18e: frame@f6e6b000(R )
  0x18f: frame@f6e6a000(R )
  0x190: frame@f6e69000(R )
  0x191: frame@f6e68000(R )
  0x192: frame@f6e67000(R )
  0x193: frame@f6e66000(R )
  0x194: frame@f6e65000(R )
  0x195: frame@f6e64000(R )
  0x196: frame@f6e63000(R )
  0x197: frame@f6e62000(R )
  0x198: frame@f6e61000(R )
  0x199: frame@f6e60000(R )
  0x19a: frame@f6e5f000(R )
  0x19b: frame@f6e5e000(R )
  0x19c: frame@f6e5d000(R )
  0x19d: frame@f6e5c000(R )
  0x19e: frame@f6e5b000(R )
  0x19f: frame@f6e5a000(R )
  0x1a0: frame@f6e59000(R )
  0x1a1: frame@f6e58000(R )
  0x1a2: frame@f6e57000(R )
  0x1a3: frame@f6e56000(R )
  0x1a4: frame@f6e55000(R )
  0x1a5: frame@f6e54000(R )
  0x1a6: frame@f6e53000(R )
  0x1a7: frame@f6e52000(R )
  0x1a8: frame@f6e51000(R )
  0x1a9: frame@f6e50000(R )
  0x1aa: frame@f6e4f000(R )
  0x1ab: frame@f6e4e000(R )
  0x1ac: frame@f6e4d000(R )
  0x1ad: frame@f6e4c000(R )
  0x1ae: frame@f6e4b000(R )
  0x1af: frame@f6e4a000(R )
  0x1b0: frame@f6e49000(R )
  0x1b1: frame@f6e48000(R )
  0x1b2: frame@f6e47000(R )
  0x1b3: frame@f6e46000(R )
  0x1b4: frame@f6e45000(R )
  0x1b5: frame@f6e44000(R )
  0x1b6: frame@f6e43000(R )
  0x1b7: frame@f6e42000(R )
  0x1b8: frame@f6e41000(R )
  0x1b9: frame@f6e40000(R )
  0x1ba: frame@f6e3f000(R )
  0x1bb: frame@f6e3e000(R )
  0x1bc: frame@f6e3d000(R )
  0x1bd: frame@f6e3c000(R )
  0x1be: frame@f6e3b000(R )
  0x1bf: frame@f6e3a000(R )
  0x1c0: frame@f6e39000(R )
  0x1c1: frame@f6e38000(R )
  0x1c2: frame@f6e37000(R )
  0x1c3: frame@f6e36000(R )
  0x1c4: frame@f6e35000(R )
  0x1c5: frame@f6e34000(R )
  0x1c6: frame@f6e33000(R )
  0x1c7: frame@f6e32000(R )
  0x1c8: frame@f6e31000(R )
  0x1c9: frame@f6e30000(R )
  0x1ca: frame@f6e2f000(R )
  0x1cb: frame@f6e2e000(R )
  0x1cc: frame@f6e2d000(R )
  0x1cd: frame@f6e2c000(R )
  0x1ce: frame@f6e2b000(R )
  0x1cf: frame@f6e2a000(R )
  0x1d0: frame@f6e29000(R )
  0x1d1: frame@f6e28000(R )
  0x1d2: frame@f6e27000(R )
  0x1d3: frame@f6e26000(R )
  0x1d4: frame@f6e25000(R )
  0x1d5: frame@f6e24000(R )
  0x1d6: frame@f6e23000(R )
  0x1d7: frame@f6e22000(R )
  0x1d8: frame@f6e21000(R )
  0x1d9: frame@f6e20000(R )
  0x1da: frame@f6e1f000(R )
  0x1db: frame@f6e1e000(R )
  0x1dc: frame@f6e1d000(R )
  0x1dd: frame@f6e1c000(R )
  0x1de: frame@f6e1b000(R )
  0x1df: frame@f6e1a000(R )
  0x1e0: frame@f6e19000(R )
  0x1e1: frame@f6e18000(R )
  0x1e2: frame@f6e17000(R )
  0x1e3: frame@f6e16000(R )
  0x1e4: frame@f6e15000(R )
  0x1e5: frame@f6e14000(R )
  0x1e6: frame@f6e13000(R )
  0x1e7: frame@f6e12000(R )
  0x1e8: frame@f6e11000(R )
  0x1e9: frame@f6e10000(R )
  0x1ea: frame@f6e0f000(R )
  0x1eb: frame@f6e0e000(R )
  0x1ec: frame@f6e0d000(R )
  0x1ed: frame@f6e0c000(R )
  0x1ee: frame@f6e0b000(R )
  0x1ef: frame@f6e0a000(R )
  0x1f0: frame@f6e09000(R )
  0x1f1: frame@f6e08000(R )
  0x1f2: frame@f6e07000(R )
  0x1f3: frame@f6e06000(R )
  0x1f4: frame@f6e05000(R )
  0x1f5: frame@f6e04000(R )
  0x1f6: frame@f6e03000(R )
  0x1f7: frame@f6e02000(R )
  0x1f8: frame@f6e01000(R )
  0x1f9: frame@f6e00000(R )
  0x1fa: frame@f6fff000(R )
  0x1fb: frame@f6ffe000(R )
  0x1fc: frame@f6ffd000(R )
  0x1fd: frame@f6ffc000(R )
  0x1fe: frame@f6ffb000(R )
  0x1ff: frame@f6ffa000(R )
  0x200: frame@f6ff9000(R )
  0x201: frame@f6ff8000(R )
  0x202: frame@f6ff7000(R )
  0x203: frame@f6ff6000(R )
  0x204: frame@f6ff5000(R )
  0x205: frame@f6ff4000(R )
  0x206: frame@f6ff3000(R )
  0x207: frame@f6ff2000(R )
  0x208: frame@f6ff1000(R )
  0x209: frame@f6ff0000(R )
  0x20a: frame@f6fef000(R )
  0x20b: frame@f6fee000(R )
  0x20c: frame@f6fed000(R )
  0x20d: frame@f6fec000(R )
  0x20e: frame@f6feb000(R )
  0x20f: frame@f6fea000(R )
  0x210: frame@f6fe9000(R )
  0x211: frame@f6fe8000(R )
  0x212: frame@f6fe7000(R )
  0x213: frame@f6fe6000(R )
  0x214: frame@f6fe5000(R )
  0x215: frame@f6fe4000(R )
  0x216: frame@f6fe3000(R )
  0x217: frame@f6fe2000(R )
  0x218: frame@f6fe1000(R )
  0x219: frame@f6fe0000(R )
  0x21a: frame@f6fdf000(R )
  0x21b: frame@f6fde000(R )
  0x21c: frame@f6fdd000(R )
  0x21d: frame@f6fdc000(R )
  0x21e: frame@f6fdb000(R )
  0x21f: frame@f6fda000(R )
  0x220: frame@f6fd9000(R )
  0x221: frame@f6fd8000(R )
  0x222: frame@f6fd7000(R )
  0x223: frame@f6fd6000(R )
  0x224: frame@f6fd5000(R )
  0x225: frame@f6fd4000(R )
  0x226: frame@f6fd3000(R )
  0x227: frame@f6fd2000(R )
  0x228: frame@f6fd1000(R )
  0x229: frame@f6fd0000(R )
  0x22a: frame@f6fcf000(R )
  0x22b: frame@f6fce000(R )
  0x22c: frame@f6fcd000(R )
  0x22d: frame@f6fcc000(R )
  0x22e: frame@f6fcb000(R )
  0x22f: frame@f6fca000(R )
  0x230: frame@f6fc9000(R )
  0x231: frame@f6fc8000(R )
  0x232: frame@f6fc7000(R )
  0x233: frame@f6fc6000(R )
  0x234: frame@f6fc5000(R )
  0x235: frame@f6fc4000(R )
  0x236: frame@f6fc3000(R )
  0x237: frame@f6fc2000(R )
  0x238: frame@f6fc1000(R )
  0x239: frame@f6fc0000(R )
  0x23a: frame@f6fbf000(R )
  0x23b: frame@f6fbe000(R )
  0x23c: frame@f6fbd000(R )
  0x23d: frame@f6fbc000(R )
  0x23e: frame@f6fbb000(R )
  0x23f: frame@f6fba000(R )
  0x240: frame@f6fb9000(R )
  0x241: frame@f6fb8000(R )
  0x242: frame@f6fb7000(R )
  0x243: frame@f6fb6000(R )
  0x244: frame@f6fb5000(R )
  0x245: frame@f6fb4000(R )
  0x246: frame@f6fb3000(R )
  0x247: frame@f6fb2000(R )
  0x248: frame@f6fb1000(R )
  0x249: frame@f6fb0000(R )
  0x24a: frame@f6faf000(R )
  0x24b: frame@f6fae000(R )
  0x24c: frame@f6fad000(R )
  0x24d: frame@f6fac000(R )
  0x24e: frame@f6fab000(R )
  0x24f: frame@f6faa000(R )
  0x250: frame@f6fa9000(R )
  0x251: frame@f6fa8000(R )
  0x252: frame@f6fa7000(R )
  0x253: frame@f6fa6000(R )
  0x254: frame@f6fa5000(R )
  0x255: frame@f6fa4000(R )
  0x256: frame@f6fa3000(R )
  0x257: frame@f6fa2000(R )
  0x258: frame@f6fa1000(R )
  0x259: frame@f6fa0000(R )
  0x25a: frame@f6f9f000(R )
  0x25b: frame@f6f9e000(R )
  0x25c: frame@f6f9d000(R )
  0x25d: frame@f6f9c000(R )
  0x25e: frame@f6f9b000(R )
  0x25f: frame@f6f9a000(R )
  0x260: frame@f6f99000(R )
  0x261: frame@f6f98000(R )
  0x262: frame@f6f97000(R )
  0x263: frame@f6f96000(R )
  0x264: frame@f6f95000(R )
  0x265: frame@f6f94000(R )
  0x266: frame@f6f93000(R )
  0x267: frame@f6f92000(R )
  0x268: frame@f6f91000(R )
  0x269: frame@f6f90000(R )
  0x26a: frame@f6f8f000(R )
  0x26b: frame@f6f8e000(R )
  0x26c: frame@f6f8d000(R )
  0x26d: frame@f6f8c000(R )
  0x26e: frame@f6f8b000(R )
  0x26f: frame@f6f8a000(R )
  0x270: frame@f6f89000(R )
  0x271: frame@f6f88000(R )
  0x272: frame@f6f87000(R )
  0x273: frame@f6f86000(R )
  0x274: frame@f6f85000(R )
  0x275: frame@f6f84000(R )
  0x276: frame@f6f83000(R )
  0x277: frame@f6f82000(R )
  0x278: frame@f6f81000(R )
  0x279: frame@f6f80000(R )
  0x27a: frame@f6f7f000(R )
  0x27b: frame@f6f7e000(R )
  0x27c: frame@f6f7d000(R )
  0x27d: frame@f6f7c000(R )
  0x27e: frame@f6f7b000(R )
  0x27f: frame@f6f7a000(R )
  0x280: frame@f6f79000(R )
  0x281: frame@f6f78000(R )
  0x282: frame@f6f77000(R )
  0x283: frame@f6f76000(R )
  0x284: frame@f6f75000(R )
  0x285: frame@f6f74000(R )
  0x286: frame@f6f73000(R )
  0x287: frame@f6f72000(R )
  0x288: frame@f6f71000(R )
  0x289: frame@f6f70000(R )
  0x28a: frame@f6f6f000(R )
  0x28b: frame@f6f6e000(R )
  0x28c: frame@f6f6d000(R )
  0x28d: frame@f6f6c000(R )
  0x28e: frame@f6f6b000(R )
  0x28f: frame@f6f6a000(R )
  0x290: frame@f6f69000(R )
  0x291: frame@f6f68000(R )
  0x292: frame@f6f67000(R )
  0x293: frame@f6f66000(R )
  0x294: frame@f6f65000(R )
  0x295: frame@f6f64000(R )
  0x296: frame@f6f63000(R )
  0x297: frame@f6f62000(R )
  0x298: frame@f6f61000(R )
  0x299: frame@f6f60000(R )
  0x29a: frame@f6f5f000(R )
  0x29b: frame@f6f5e000(R )
  0x29c: frame@f6f5d000(R )
  0x29d: frame@f6f5c000(R )
  0x29e: frame@f6f5b000(R )
  0x29f: frame@f6f5a000(R )
  0x2a0: frame@f6f59000(R )
  0x2a1: frame@f6f58000(R )
  0x2a2: frame@f6f57000(R )
  0x2a3: frame@f6f56000(R )
  0x2a4: frame@f6f55000(R )
  0x2a5: frame@f6f54000(R )
  0x2a6: frame@f6f53000(R )
  0x2a7: frame@f6f52000(R )
  0x2a8: frame@f6f51000(R )
  0x2a9: frame@f6f50000(R )
  0x2aa: frame@f6f4f000(R )
  0x2ab: frame@f6f4e000(R )
  0x2ac: frame@f6f4d000(R )
  0x2ad: frame@f6f4c000(R )
  0x2ae: frame@f6f4b000(R )
  0x2af: frame@f6f4a000(R )
  0x2b0: frame@f6f49000(R )
  0x2b1: frame@f6f48000(R )
  0x2b2: frame@f6f47000(R )
  0x2b3: frame@f6f46000(R )
  0x2b4: frame@f6f45000(R )
  0x2b5: frame@f6f44000(R )
  0x2b6: frame@f6f43000(R )
  0x2b7: frame@f6f42000(R )
  0x2b8: frame@f6f41000(R )
  0x2b9: frame@f6f40000(R )
  0x2ba: frame@f6f3f000(R )
  0x2bb: frame@f6f3e000(R )
  0x2bc: frame@f6f3d000(R )
  0x2bd: frame@f6f3c000(R )
  0x2be: frame@f6f3b000(R )
  0x2bf: frame@f6f3a000(R )
  0x2c0: frame@f6f39000(R )
  0x2c1: frame@f6f38000(R )
  0x2c2: frame@f6f37000(R )
  0x2c3: frame@f6f36000(R )
  0x2c4: frame@f6f35000(R )
  0x2c5: frame@f6f34000(R )
  0x2c6: frame@f6f33000(R )
  0x2c7: frame@f6f32000(R )
  0x2c8: frame@f6f31000(R )
  0x2c9: frame@f6f30000(R )
  0x2ca: frame@f6f2f000(R )
  0x2cb: frame@f6f2e000(R )
  0x2cc: frame@f6f2d000(R )
  0x2cd: frame@f6f2c000(R )
  0x2ce: frame@f6f2b000(R )
  0x2cf: frame@f6f2a000(R )
  0x2d0: frame@f6f29000(R )
  0x2d1: frame@f6f28000(R )
  0x2d2: frame@f6f27000(R )
  0x2d3: frame@f6f26000(R )
  0x2d4: frame@f6f25000(R )
  0x2d5: frame@f6f24000(R )
  0x2d6: frame@f6f23000(R )
  0x2d7: frame@f6f22000(R )
  0x2d8: frame@f6f21000(R )
  0x2d9: frame@f6f20000(R )
  0x2da: frame@f6f1f000(R )
  0x2db: frame@f6f1e000(R )
  0x2dc: frame@f6f1d000(R )
  0x2dd: frame@f6f1c000(R )
  0x2de: frame@f6f1b000(R )
  0x2df: frame@f6f1a000(R )
  0x2e0: frame@f6f19000(R )
  0x2e1: frame@f6f18000(R )
  0x2e2: frame@f6f17000(R )
  0x2e3: frame@f6f16000(R )
  0x2e4: frame@f6f15000(R )
  0x2e5: frame@f6f14000(R )
  0x2e6: frame@f6f13000(R )
  0x2e7: frame@f6f12000(R )
  0x2e8: frame@f6f11000(R )
  0x2e9: frame@f6f10000(R )
  0x2ea: frame@f6f0f000(R )
  0x2eb: frame@f6f0e000(R )
  0x2ec: frame@f6f0d000(R )
  0x2ed: frame@f6f0c000(R )
  0x2ee: frame@f6f0b000(R )
  0x2ef: frame@f6f0a000(R )
  0x2f0: frame@f6f09000(R )
  0x2f1: frame@f6f08000(R )
  0x2f2: frame@f6f07000(R )
  0x2f3: frame@f6f06000(R )
  0x2f4: frame@f6f05000(R )
  0x2f5: frame@f6f04000(R )
  0x2f6: frame@f6f03000(R )
  0x2f7: frame@f6f02000(R )
  0x2f8: frame@f6f01000(R )
  0x2f9: frame@f6f00000(R )
  0x2fa: frame@f70ff000(R )
  0x2fb: frame@f70fe000(R )
  0x2fc: frame@f70fd000(R )
  0x2fd: frame@f70fc000(R )
  0x2fe: frame@f70fb000(R )
  0x2ff: frame@f70fa000(R )
  0x300: frame@f70f9000(R )
  0x301: frame@f70f8000(R )
  0x302: frame@f70f7000(R )
  0x303: frame@f70f6000(R )
  0x304: frame@f70f5000(R )
  0x305: frame@f70f4000(R )
  0x306: frame@f70f3000(R )
  0x307: frame@f70f2000(R )
  0x308: frame@f70f1000(R )
  0x309: frame@f70f0000(R )
  0x30a: frame@f70ef000(R )
  0x30b: frame@f70ee000(R )
  0x30c: frame@f70ed000(R )
  0x30d: frame@f70ec000(R )
  0x30e: frame@f70eb000(R )
  0x30f: frame@f70ea000(R )
  0x310: frame@f70e9000(R )
  0x311: frame@f70e8000(R )
  0x312: frame@f70e7000(R )
  0x313: frame@f70e6000(R )
  0x314: frame@f70e5000(R )
  0x315: frame@f70e4000(R )
  0x316: frame@f70e3000(R )
  0x317: frame@f70e2000(R )
  0x318: frame@f70e1000(R )
  0x319: frame@f70e0000(R )
  0x31a: frame@f70df000(R )
  0x31b: frame@f70de000(R )
  0x31c: frame@f70dd000(R )
  0x31d: frame@f70dc000(R )
  0x31e: frame@f70db000(R )
  0x31f: frame@f70da000(R )
  0x320: frame@f70d9000(R )
  0x321: frame@f70d8000(R )
  0x322: frame@f70d7000(R )
  0x323: frame@f70d6000(R )
  0x324: frame@f70d5000(R )
  0x325: frame@f70d4000(R )
  0x326: frame@f70d3000(R )
  0x327: frame@f70d2000(R )

  0x328: frame@f70d1000(R )
  0x329: frame@f70d0000(R )
  0x32a: frame@f70cf000(R )
  0x32b: frame@f70ce000(R )
  0x32c: frame@f70cd000(R )
  0x32d: frame@f70cc000(R )
  0x32e: frame@f70cb000(R )
  0x32f: frame@f70ca000(R )
  0x330: frame@f70c9000(R )
  0x331: frame@f70c8000(R )
  0x332: frame@f70c7000(R )
  0x333: frame@f70c6000(R )
  0x334: frame@f70c5000(R )
  0x335: frame@f70c4000(R )
  0x336: frame@f70c3000(R )
  0x337: frame@f70c2000(R )
  0x338: frame@f70c1000(R )
  0x339: frame@f70c0000(R )
  0x33a: frame@f70bf000(R )
  0x33b: frame@f70be000(R )
  0x33c: frame@f70bd000(R )
  0x33d: frame@f70bc000(R )
  0x33e: frame@f70bb000(R )
  0x33f: frame@f70ba000(R )
  0x340: frame@f70b9000(R )
  0x341: frame@f70b8000(R )
  0x342: frame@f70b7000(R )
  0x343: frame@f70b6000(R )
  0x344: frame@f70b5000(R )
  0x345: frame@f70b4000(R )
  0x346: frame@f70b3000(R )
  0x347: frame@f70b2000(R )
  0x348: frame@f70b1000(R )
  0x349: frame@f70b0000(R )
  0x34a: frame@f70af000(R )
  0x34b: frame@f70ae000(R )
  0x34c: frame@f70ad000(R )
  0x34d: frame@f70ac000(R )
  0x34e: frame@f70ab000(R )
  0x34f: frame@f70aa000(R )
  0x350: frame@f70a9000(R )
  0x351: frame@f70a8000(R )
  0x352: frame@f70a7000(R )
  0x353: frame@f70a6000(R )
  0x354: frame@f70a5000(R )
  0x355: frame@f70a4000(R )
  0x356: frame@f70a3000(R )
  0x357: frame@f70a2000(R )
  0x358: frame@f70a1000(R )
  0x359: frame@f70a0000(R )
  0x35a: frame@f709f000(R )
  0x35b: frame@f709e000(R )
  0x35c: frame@f709d000(R )
  0x35d: frame@f709c000(R )
  0x35e: frame@f709b000(R )
  0x35f: frame@f709a000(R )
  0x360: frame@f7099000(R )
  0x361: frame@f7098000(R )
  0x362: frame@f7097000(R )
  0x363: frame@f7096000(R )
  0x364: frame@f7095000(R )
  0x365: frame@f7094000(R )
  0x366: frame@f7093000(R )
  0x367: frame@f7092000(R )
  0x368: frame@f7091000(R )
  0x369: frame@f7090000(R )
  0x36a: frame@f708f000(R )
  0x36b: frame@f708e000(R )
  0x36c: frame@f708d000(R )
  0x36d: frame@f708c000(R )
  0x36e: frame@f708b000(R )
  0x36f: frame@f708a000(R )
  0x370: frame@f7089000(R )
  0x371: frame@f7088000(R )
  0x372: frame@f7087000(R )
  0x373: frame@f7086000(R )
  0x374: frame@f7085000(R )
  0x375: frame@f7084000(R )
  0x376: frame@f7083000(R )
  0x377: frame@f7082000(R )
  0x378: frame@f7081000(R )
  0x379: frame@f7080000(R )
  0x37a: frame@f707f000(R )
  0x37b: frame@f707e000(R )
  0x37c: frame@f707d000(R )
  0x37d: frame@f707c000(R )
  0x37e: frame@f707b000(R )
  0x37f: frame@f707a000(R )
  0x380: frame@f7079000(R )
  0x381: frame@f7078000(R )
  0x382: frame@f7077000(R )
  0x383: frame@f7076000(R )
  0x384: frame@f7075000(R )
  0x385: frame@f7074000(R )
  0x386: frame@f7073000(R )
  0x387: frame@f7072000(R )
  0x388: frame@f7071000(R )
  0x389: frame@f7070000(R )
  0x38a: frame@f706f000(R )
  0x38b: frame@f706e000(R )
  0x38c: frame@f706d000(R )
  0x38d: frame@f706c000(R )
  0x38e: frame@f706b000(R )
  0x38f: frame@f706a000(R )
  0x390: frame@f7069000(R )
  0x391: frame@f7068000(R )
  0x392: frame@f7067000(R )
  0x393: frame@f7066000(R )
  0x394: frame@f7065000(R )
  0x395: frame@f7064000(R )
  0x396: frame@f7063000(R )
  0x397: frame@f7062000(R )
  0x398: frame@f7061000(R )
  0x399: frame@f7060000(R )
  0x39a: frame@f705f000(R )
  0x39b: frame@f705e000(R )
  0x39c: frame@f705d000(R )
  0x39d: frame@f705c000(R )
  0x39e: frame@f705b000(R )
  0x39f: frame@f705a000(R )
  0x3a0: frame@f7059000(R )
  0x3a1: frame@f7058000(R )
  0x3a2: frame@f7057000(R )
  0x3a3: frame@f7056000(R )
  0x3a4: frame@f7055000(R )
  0x3a5: frame@f7054000(R )
  0x3a6: frame@f7053000(R )
  0x3a7: frame@f7052000(R )
  0x3a8: frame@f7051000(R )
  0x3a9: frame@f7050000(R )
  0x3aa: frame@f704f000(R )
  0x3ab: frame@f704e000(R )
  0x3ac: frame@f704d000(R )
  0x3ad: frame@f704c000(R )
  0x3ae: frame@f704b000(R )
  0x3af: frame@f704a000(R )
  0x3b0: frame@f7049000(R )
  0x3b1: frame@f7048000(R )
  0x3b2: frame@f7047000(R )
  0x3b3: frame@f7046000(R )
  0x3b4: frame@f7045000(R )
  0x3b5: frame@f7044000(R )
  0x3b6: frame@f7043000(R )
  0x3b7: frame@f7042000(R )
  0x3b8: frame@f7041000(R )
  0x3b9: frame@f7040000(R )
  0x3ba: frame@f703f000(R )
  0x3bb: frame@f703e000(R )
  0x3bc: frame@f703d000(R )
  0x3bd: frame@f703c000(R )
  0x3be: frame@f703b000(R )
  0x3bf: frame@f703a000(R )
  0x3c0: frame@f7039000(R )
  0x3c1: frame@f7038000(R )
  0x3c2: frame@f7037000(R )
  0x3c3: frame@f7036000(R )
  0x3c4: frame@f7035000(R )
  0x3c5: frame@f7034000(R )
  0x3c6: frame@f7033000(R )
  0x3c7: frame@f7032000(R )
  0x3c8: frame@f7031000(R )
  0x3c9: frame@f7030000(R )
  0x3ca: frame@f702f000(R )
  0x3cb: frame@f702e000(R )
  0x3cc: frame@f702d000(R )
  0x3cd: frame@f702c000(R )
  0x3ce: frame@f702b000(R )
  0x3cf: frame@f702a000(R )
  0x3d0: frame@f7029000(R )
  0x3d1: frame@f7028000(R )
  0x3d2: frame@f7027000(R )
  0x3d3: frame@f7026000(R )
  0x3d4: frame@f7025000(R )
  0x3d5: frame@f7024000(R )
  0x3d6: frame@f7023000(R )
  0x3d7: frame@f7022000(R )
  0x3d8: frame@f7021000(R )
  0x3d9: frame@f7020000(R )
  0x3da: frame@f701f000(R )
  0x3db: frame@f701e000(R )
  0x3dc: frame@f701d000(R )
  0x3dd: frame@f701c000(R )
  0x3de: frame@f701b000(R )
  0x3df: frame@f701a000(R )
  0x3e0: frame@f7019000(R )
  0x3e1: frame@f7018000(R )
  0x3e2: frame@f7017000(R )
  0x3e3: frame@f7016000(R )
  0x3e4: frame@f7015000(R )
  0x3e5: frame@f7014000(R )
  0x3e6: frame@f7013000(R )
  0x3e7: frame@f7012000(R )
  0x3e8: frame@f7011000(R )
  0x3e9: frame@f7010000(R )
  0x3ea: frame@f700f000(R )
  0x3eb: frame@f700e000(R )
  0x3ec: frame@f700d000(R )
  0x3ed: frame@f700c000(R )
  0x3ee: frame@f700b000(R )
  0x3ef: frame@f700a000(R )
  0x3f0: frame@f7009000(R )
  0x3f1: frame@f7008000(R )
  0x3f2: frame@f7007000(R )
  0x3f3: frame@f7006000(R )
  0x3f4: frame@f7005000(R )
  0x3f5: frame@f7004000(R )
  0x3f6: frame@f7003000(R )
  0x3f7: frame@f7002000(R )
  0x3f8: frame@f7001000(R )
  0x3f9: frame@f7000000(R )
  0x3fa: frame@f71ff000(R )
  0x3fb: frame@f71fe000(R )
  0x3fc: frame@f71fd000(R )
  0x3fd: frame@f71fc000(R )
  0x3fe: frame@f71fb000(R )
  0x3ff: frame@f71fa000(R )
}
pt@f6df3000{
  0x0: frame@f729d000(RW)
  0x1: frame@f9dc2000(RW)
  0x2: frame@f9dc3000(RW)
}
pt@f6df6000{
  0x180: frame@d0180000(RW)
  0x181: frame@d0181000(RW)
  0x182: frame@d0182000(RW)
  0x183: frame@d0183000(RW)
  0x184: frame@d0184000(RW)
  0x185: frame@d0185000(RW)
  0x186: frame@d0186000(RW)
  0x187: frame@d0187000(RW)
  0x188: frame@d0188000(RW)
  0x189: frame@d0189000(RW)
  0x18a: frame@d018a000(RW)
  0x18b: frame@d018b000(RW)
  0x18c: frame@d018c000(RW)
  0x18d: frame@d018d000(RW)
  0x18e: frame@d018e000(RW)
  0x18f: frame@d018f000(RW)
  0x190: frame@d0190000(RW)
  0x191: frame@d0191000(RW)
  0x192: frame@d0192000(RW)
  0x193: frame@d0193000(RW)
  0x194: frame@d0194000(RW)
  0x195: frame@d0195000(RW)
  0x196: frame@d0196000(RW)
  0x197: frame@d0197000(RW)
  0x198: frame@d0198000(RW)
  0x199: frame@d0199000(RW)
  0x19a: frame@d019a000(RW)
  0x19b: frame@d019b000(RW)
  0x19c: frame@d019c000(RW)
  0x19d: frame@d019d000(RW)
  0x19e: frame@d019e000(RW)
  0x19f: frame@d019f000(RW)
  0x1a5: frame@d01a5000(RW)
}
pt@f6df7000{
  0x0: frame@f9a6c000(RW)
  0x1: frame@f9a6b000(RW)
  0x2: frame@f9a6a000(RW)
  0x3: frame@f9a69000(RW)
  0x4: frame@f9a68000(RW)
  0x5: frame@f9a67000(RW)
  0x6: frame@f9a66000(RW)
  0x7: frame@f9a65000(RW)
  0x8: frame@f9a64000(RW)
  0x9: frame@f9a63000(RW)
  0xa: frame@f9a62000(RW)
  0xb: frame@f9a61000(RW)
  0xc: frame@f9a60000(RW)
  0xd: frame@f9a5f000(RW)
  0xe: frame@f9a5e000(RW)
  0xf: frame@f9a5d000(RW)
  0x10: frame@f9a5c000(RW)
  0x11: frame@f9a5b000(RW)
  0x12: frame@f9a5a000(RW)
  0x13: frame@f9a59000(RW)
  0x14: frame@f9a58000(RW)
  0x15: frame@f9a57000(RW)
  0x16: frame@f9a56000(RW)
  0x17: frame@f9a55000(RW)
  0x18: frame@f9a54000(RW)
  0x19: frame@f9a53000(RW)
  0x1a: frame@f9a52000(RW)
  0x1b: frame@f9a51000(RW)
  0x1c: frame@f9a50000(RW)
  0x1d: frame@f9a4f000(RW)
  0x1e: frame@f9a4e000(RW)
  0x1f: frame@f9a4d000(RW)
  0x20: frame@f9a4c000(RW)
  0x21: frame@f9a4b000(RW)
  0x22: frame@f9a4a000(RW)
  0x23: frame@f9a49000(RW)
  0x24: frame@f9a48000(RW)
  0x25: frame@f9a47000(RW)
  0x26: frame@f9a46000(RW)
  0x27: frame@f9a45000(RW)
  0x28: frame@f9a44000(RW)
  0x29: frame@f9a43000(RW)
  0x2a: frame@f9a42000(RW)
  0x2b: frame@f9a41000(RW)
  0x2c: frame@f9a40000(RW)
  0x2d: frame@f9a3f000(RW)
  0x2e: frame@f9a3e000(RW)
  0x2f: frame@f9a3d000(RW)
  0x30: frame@f9a3c000(RW)
  0x31: frame@f9a3b000(RW)
  0x32: frame@f9a3a000(RW)
  0x33: frame@f9a39000(RW)
  0x34: frame@f9a38000(RW)
  0x35: frame@f9a37000(RW)
  0x36: frame@f9a36000(RW)
  0x37: frame@f9a35000(RW)
  0x38: frame@f9a34000(RW)
  0x39: frame@f9a33000(RW)
  0x3a: frame@f9a32000(RW)
  0x3b: frame@f9a31000(RW)
  0x3c: frame@f9a30000(RW)
  0x3d: frame@f9a2f000(RW)
  0x3e: frame@f9a2e000(RW)
  0x3f: frame@f9a2d000(RW)
  0x40: frame@f9a2c000(RW)
  0x41: frame@f9a2b000(RW)
  0x42: frame@f9a2a000(RW)
  0x43: frame@f9a29000(RW)
  0x44: frame@f9a28000(RW)
  0x45: frame@f9a27000(RW)
  0x46: frame@f9a26000(RW)
  0x47: frame@f9a25000(RW)
  0x48: frame@f9a24000(RW)
  0x49: frame@f9a23000(RW)
  0x4a: frame@f9a22000(RW)
  0x4b: frame@f9a21000(RW)
  0x4c: frame@f9a20000(RW)
  0x4d: frame@f9a1f000(RW)
  0x4e: frame@f9a1e000(RW)
  0x4f: frame@f9a1d000(RW)
  0x50: frame@f9a1c000(RW)
  0x51: frame@f9a1b000(RW)
  0x52: frame@f9a1a000(RW)
  0x53: frame@f9a19000(RW)
  0x54: frame@f9a18000(RW)
  0x55: frame@f9a17000(RW)
  0x56: frame@f9a16000(RW)
  0x57: frame@f9a15000(RW)
  0x58: frame@f9a14000(RW)
  0x59: frame@f9a13000(RW)
  0x5a: frame@f9a12000(RW)
  0x5b: frame@f9a11000(RW)
  0x5c: frame@f9a10000(RW)
  0x5d: frame@f9a0f000(RW)
  0x5e: frame@f9a0e000(RW)
  0x5f: frame@f9a0d000(RW)
  0x60: frame@f9a0c000(RW)
  0x61: frame@f9a0b000(RW)
  0x62: frame@f9a0a000(RW)
  0x63: frame@f9a09000(RW)
  0x64: frame@f9a08000(RW)
  0x65: frame@f9a07000(RW)
  0x66: frame@f9a06000(RW)
  0x67: frame@f9a05000(RW)
  0x68: frame@f9a04000(RW)
  0x69: frame@f9a03000(RW)
  0x6a: frame@f9a02000(RW)
  0x6b: frame@f9a01000(RW)
  0x6c: frame@f9a00000(RW)
  0x6d: frame@f9bff000(RW)
  0x6e: frame@f9bfe000(RW)
  0x6f: frame@f9bfd000(RW)
  0x70: frame@f9bfc000(RW)
  0x71: frame@f9bfb000(RW)
  0x72: frame@f9bfa000(RW)
  0x73: frame@f9bf9000(RW)
  0x74: frame@f9bf8000(RW)
  0x75: frame@f9bf7000(RW)
  0x76: frame@f9bf6000(RW)
  0x77: frame@f9bf5000(RW)
  0x78: frame@f9bf4000(RW)
  0x79: frame@f9bf3000(RW)
  0x7a: frame@f9bf2000(RW)
  0x7b: frame@f9bf1000(RW)
  0x7c: frame@f9bf0000(RW)
  0x7d: frame@f9bef000(RW)
  0x7e: frame@f9bee000(RW)
  0x7f: frame@f9bed000(RW)
  0x80: frame@f9bec000(RW)
  0x81: frame@f9beb000(RW)
  0x82: frame@f9bea000(RW)
  0x83: frame@f9be9000(RW)
  0x84: frame@f9be8000(RW)
  0x85: frame@f9be7000(RW)
  0x86: frame@f9be6000(RW)
  0x87: frame@f9be5000(RW)
  0x88: frame@f9be4000(RW)
  0x89: frame@f9be3000(RW)
  0x8a: frame@f9be2000(RW)
  0x8b: frame@f9be1000(RW)
  0x8c: frame@f9be0000(RW)
  0x8d: frame@f9bdf000(RW)
  0x8e: frame@f9bde000(RW)
  0x8f: frame@f9bdd000(RW)
  0x90: frame@f9bdc000(RW)
  0x91: frame@f9bdb000(RW)
  0x92: frame@f9bda000(RW)
  0x93: frame@f9bd9000(RW)
  0x94: frame@f9bd8000(RW)
  0x95: frame@f9bd7000(RW)
  0x96: frame@f9bd6000(RW)
  0x97: frame@f9bd5000(RW)
  0x98: frame@f9bd4000(RW)
  0x99: frame@f9bd3000(RW)
  0x9a: frame@f9bd2000(RW)
  0x9b: frame@f9bd1000(RW)
  0x9c: frame@f9bd0000(RW)
  0x9d: frame@f9bcf000(RW)
  0x9e: frame@f9bce000(RW)
  0x9f: frame@f9bcd000(RW)
  0xa0: frame@f9bcc000(RW)
  0xa1: frame@f9bcb000(RW)
  0xa2: frame@f9bca000(RW)
  0xa3: frame@f9bc9000(RW)
  0xa4: frame@f9bc8000(RW)
  0xa5: frame@f9bc7000(RW)
  0xa6: frame@f9bc6000(RW)
  0xa7: frame@f9bc5000(RW)
  0xa8: frame@f9bc4000(RW)
  0xa9: frame@f9bc3000(RW)
  0xaa: frame@f9bc2000(RW)
  0xab: frame@f9bc1000(RW)
  0xac: frame@f9bc0000(RW)
  0xad: frame@f9bbf000(RW)
  0xae: frame@f9bbe000(RW)
  0xaf: frame@f9bbd000(RW)
  0xb0: frame@f9bbc000(RW)
  0xb1: frame@f9bbb000(RW)
  0xb2: frame@f9bba000(RW)
  0xb3: frame@f9bb9000(RW)
  0xb4: frame@f9bb8000(RW)
  0xb5: frame@f9bb7000(RW)
  0xb6: frame@f9bb6000(RW)
  0xb7: frame@f9bb5000(RW)
  0xb8: frame@f9bb4000(RW)
  0xb9: frame@f9bb3000(RW)
  0xba: frame@f9bb2000(RW)
  0xbb: frame@f9bb1000(RW)
  0xbc: frame@f9bb0000(RW)
  0xbd: frame@f9baf000(RW)
  0xbe: frame@f9bae000(RW)
  0xbf: frame@f9bad000(RW)
  0xc0: frame@f9bac000(RW)
  0xc1: frame@f9bab000(RW)
  0xc2: frame@f9baa000(RW)
  0xc3: frame@f9ba9000(RW)
  0xc4: frame@f9ba8000(RW)
  0xc5: frame@f9ba7000(RW)
  0xc6: frame@f9ba6000(RW)
  0xc7: frame@f9ba5000(RW)
  0xc8: frame@f9ba4000(RW)
  0xc9: frame@f9ba3000(RW)
  0xca: frame@f9ba2000(RW)
  0xcb: frame@f9ba1000(RW)
  0xcc: frame@f9ba0000(RW)
  0xcd: frame@f9b9f000(RW)
  0xce: frame@f9b9e000(RW)
  0xcf: frame@f9b9d000(RW)
  0xd0: frame@f9b9c000(RW)
  0xd1: frame@f9b9b000(RW)
  0xd2: frame@f9b9a000(RW)
  0xd3: frame@f9b99000(RW)
  0xd4: frame@f9b98000(RW)
  0xd5: frame@f9b97000(RW)
  0xd6: frame@f9b96000(RW)
  0xd7: frame@f9b95000(RW)
  0xd8: frame@f9b94000(RW)
  0xd9: frame@f9b93000(RW)
  0xda: frame@f9b92000(RW)
  0xdb: frame@f9b91000(RW)
  0xdc: frame@f9b90000(RW)
  0xdd: frame@f9b8f000(RW)
  0xde: frame@f9b8e000(RW)
  0xdf: frame@f9b8d000(RW)
  0xe0: frame@f9b8c000(RW)
  0xe1: frame@f9b8b000(RW)
  0xe2: frame@f9b8a000(RW)
  0xe3: frame@f9b89000(RW)
  0xe4: frame@f9b88000(RW)
  0xe5: frame@f9b87000(RW)
  0xe6: frame@f9b86000(RW)
  0xe7: frame@f9b85000(RW)
  0xe8: frame@f9b84000(RW)
  0xe9: frame@f9b83000(RW)
  0xea: frame@f9b82000(RW)
  0xeb: frame@f9b81000(RW)
  0xec: frame@f9b80000(RW)
  0xed: frame@f9b7f000(RW)
  0xee: frame@f9b7e000(RW)
  0xef: frame@f9b7d000(RW)
  0xf0: frame@f9b7c000(RW)
  0xf1: frame@f9b7b000(RW)
  0xf2: frame@f9b7a000(RW)
  0xf3: frame@f9b79000(RW)
  0xf4: frame@f9b78000(RW)
  0xf5: frame@f9b77000(RW)
  0xf6: frame@f9b76000(RW)
  0xf7: frame@f9b75000(RW)
  0xf8: frame@f9b74000(RW)
  0xf9: frame@f9b73000(RW)
  0xfa: frame@f9b72000(RW)
  0xfb: frame@f9b71000(RW)
  0xfc: frame@f9b70000(RW)
  0xfd: frame@f9b6f000(RW)
  0xfe: frame@f9b6e000(RW)
  0xff: frame@f9b6d000(RW)
  0x100: frame@f9b6c000(RW)
  0x101: frame@f9b6b000(RW)
  0x102: frame@f9b6a000(RW)
  0x103: frame@f9b69000(RW)
  0x104: frame@f9b68000(RW)
  0x105: frame@f9b67000(RW)
  0x106: frame@f9b66000(RW)
  0x107: frame@f9b65000(RW)
  0x108: frame@f9b64000(RW)
  0x109: frame@f9b63000(RW)
  0x10a: frame@f9b62000(RW)
  0x10b: frame@f9b61000(RW)
  0x10c: frame@f9b60000(RW)
  0x10d: frame@f9b5f000(RW)
  0x10e: frame@f9b5e000(RW)
  0x10f: frame@f9b5d000(RW)
  0x110: frame@f9b5c000(RW)
  0x111: frame@f9b5b000(RW)
  0x112: frame@f9b5a000(RW)
  0x113: frame@f9b59000(RW)
  0x114: frame@f9b58000(RW)
  0x115: frame@f9b57000(RW)
  0x116: frame@f9b56000(RW)
  0x117: frame@f9b55000(RW)
  0x118: frame@f9b54000(RW)
  0x119: frame@f9b53000(RW)
  0x11a: frame@f9b52000(RW)
  0x11b: frame@f9b51000(RW)
  0x11c: frame@f9b50000(RW)
  0x11d: frame@f9b4f000(RW)
  0x11e: frame@f9b4e000(RW)
  0x11f: frame@f9b4d000(RW)
  0x120: frame@f9b4c000(RW)
  0x121: frame@f9b4b000(RW)
  0x122: frame@f9b4a000(RW)
  0x123: frame@f9b49000(RW)
  0x124: frame@f9b48000(RW)
  0x125: frame@f9b47000(RW)
  0x126: frame@f9b46000(RW)
  0x127: frame@f9b45000(RW)
  0x128: frame@f9b44000(RW)
  0x129: frame@f9b43000(RW)
  0x12a: frame@f9b42000(RW)
  0x12b: frame@f9b41000(RW)
  0x12c: frame@f9b40000(RW)
  0x12d: frame@f9b3f000(RW)
  0x12e: frame@f9b3e000(RW)
  0x12f: frame@f9b3d000(RW)
  0x130: frame@f9b3c000(RW)
  0x131: frame@f9b3b000(RW)
  0x132: frame@f9b3a000(RW)
  0x133: frame@f9b39000(RW)
  0x134: frame@f9b38000(RW)
  0x135: frame@f9b37000(RW)
  0x136: frame@f9b36000(RW)
  0x137: frame@f9b35000(RW)
  0x138: frame@f9b34000(RW)
  0x139: frame@f9b33000(RW)
  0x13a: frame@f9b32000(RW)
  0x13b: frame@f9b31000(RW)
  0x13c: frame@f9b30000(RW)
  0x13d: frame@f9b2f000(RW)
  0x13e: frame@f9b2e000(RW)
  0x13f: frame@f9b2d000(RW)
  0x140: frame@f9b2c000(RW)
  0x141: frame@f9b2b000(RW)
  0x142: frame@f9b2a000(RW)
  0x143: frame@f9b29000(RW)
  0x144: frame@f9b28000(RW)
  0x145: frame@f9b27000(RW)
  0x146: frame@f9b26000(RW)
  0x147: frame@f9b25000(RW)
  0x148: frame@f9b24000(RW)
  0x149: frame@f9b23000(RW)
  0x14a: frame@f9b22000(RW)
  0x14b: frame@f9b21000(RW)
  0x14c: frame@f9b20000(RW)
  0x14d: frame@f9b1f000(RW)
  0x14e: frame@f9b1e000(RW)
  0x14f: frame@f9b1d000(RW)
  0x150: frame@f9b1c000(RW)
  0x151: frame@f9b1b000(RW)
  0x152: frame@f9b1a000(RW)
  0x153: frame@f9b19000(RW)
  0x154: frame@f9b18000(RW)
  0x155: frame@f9b17000(RW)
  0x156: frame@f9b16000(RW)
  0x157: frame@f9b15000(RW)
  0x158: frame@f9b14000(RW)
  0x159: frame@f9b13000(RW)
  0x15a: frame@f9b12000(RW)
  0x15b: frame@f9b11000(RW)
  0x15c: frame@f9b10000(RW)
  0x15d: frame@f9b0f000(RW)
  0x15e: frame@f9b0e000(RW)
  0x15f: frame@f9b0d000(RW)
  0x160: frame@f9b0c000(RW)
  0x161: frame@f9b0b000(RW)
  0x162: frame@f9b0a000(RW)
  0x163: frame@f9b09000(RW)
  0x164: frame@f9b08000(RW)
  0x165: frame@f9b07000(RW)
  0x166: frame@f9b06000(RW)
  0x167: frame@f9b05000(RW)
  0x168: frame@f9b04000(RW)
  0x169: frame@f9b03000(RW)
  0x16a: frame@f9b02000(RW)
  0x16b: frame@f9b01000(RW)
  0x16c: frame@f9b00000(RW)
  0x16d: frame@f9cff000(RW)
  0x16e: frame@f9cfe000(RW)
  0x16f: frame@f9cfd000(RW)
  0x170: frame@f9cfc000(RW)
  0x171: frame@f9cfb000(RW)
  0x172: frame@f9cfa000(RW)
  0x173: frame@f9cf9000(RW)
  0x174: frame@f9cf8000(RW)
  0x175: frame@f9cf7000(RW)
  0x176: frame@f9cf6000(RW)
  0x177: frame@f9cf5000(RW)
  0x178: frame@f9cf4000(RW)
  0x179: frame@f9cf3000(RW)
  0x17a: frame@f9cf2000(RW)
  0x17b: frame@f9cf1000(RW)
  0x17c: frame@f9cf0000(RW)
  0x17d: frame@f9cef000(RW)
  0x17e: frame@f9cee000(RW)
  0x17f: frame@f9ced000(RW)
  0x180: frame@f9cec000(RW)
  0x181: frame@f9ceb000(RW)
  0x182: frame@f9cea000(RW)
  0x183: frame@f9ce9000(RW)
  0x184: frame@f9ce8000(RW)
  0x185: frame@f9ce7000(RW)
  0x186: frame@f9ce6000(RW)
  0x187: frame@f9ce5000(RW)
  0x188: frame@f9ce4000(RW)
  0x189: frame@f9ce3000(RW)
  0x18a: frame@f9ce2000(RW)
  0x18b: frame@f9ce1000(RW)
  0x18c: frame@f9ce0000(RW)
  0x18d: frame@f9cdf000(RW)
  0x18e: frame@f9cde000(RW)
  0x18f: frame@f9cdd000(RW)
  0x190: frame@f9cdc000(RW)
  0x191: frame@f9cdb000(RW)
  0x192: frame@f9cda000(RW)
  0x193: frame@f9cd9000(RW)
  0x194: frame@f9cd8000(RW)
  0x195: frame@f9cd7000(RW)
  0x196: frame@f9cd6000(RW)
  0x197: frame@f9cd5000(RW)
  0x198: frame@f9cd4000(RW)
  0x199: frame@f9cd3000(RW)
  0x19a: frame@f9cd2000(RW)
  0x19b: frame@f9cd1000(RW)
  0x19c: frame@f9cd0000(RW)
  0x19d: frame@f9ccf000(RW)
  0x19e: frame@f9cce000(RW)
  0x19f: frame@f9ccd000(RW)
  0x1a0: frame@f9ccc000(RW)
  0x1a1: frame@f9ccb000(RW)
  0x1a2: frame@f9cca000(RW)
  0x1a3: frame@f9cc9000(RW)
  0x1a4: frame@f9cc8000(RW)
  0x1a5: frame@f9cc7000(RW)
  0x1a6: frame@f9cc6000(RW)
  0x1a7: frame@f9cc5000(RW)
  0x1a8: frame@f9cc4000(RW)
  0x1a9: frame@f9cc3000(RW)
  0x1aa: frame@f9cc2000(RW)
  0x1ab: frame@f9cc1000(RW)
  0x1ac: frame@f9cc0000(RW)
  0x1ad: frame@f9cbf000(RW)
  0x1ae: frame@f9cbe000(RW)
  0x1af: frame@f9cbd000(RW)
  0x1b0: frame@f9cbc000(RW)
  0x1b1: frame@f9cbb000(RW)
  0x1b2: frame@f9cba000(RW)
  0x1b3: frame@f9cb9000(RW)
  0x1b4: frame@f9cb8000(RW)
  0x1b5: frame@f9cb7000(RW)
  0x1b6: frame@f9cb6000(RW)
  0x1b7: frame@f9cb5000(RW)
  0x1b8: frame@f9cb4000(RW)
  0x1b9: frame@f9cb3000(RW)
  0x1ba: frame@f9cb2000(RW)
  0x1bb: frame@f9cb1000(RW)
  0x1bc: frame@f9cb0000(RW)
  0x1bd: frame@f9caf000(RW)
  0x1be: frame@f9cae000(RW)
  0x1bf: frame@f9cad000(RW)
  0x1c0: frame@f9cac000(RW)
  0x1c1: frame@f9cab000(RW)
  0x1c2: frame@f9caa000(RW)
  0x1c3: frame@f9ca9000(RW)
  0x1c4: frame@f9ca8000(RW)
  0x1c5: frame@f9ca7000(RW)
  0x1c6: frame@f9ca6000(RW)
  0x1c7: frame@f9ca5000(RW)
  0x1c8: frame@f9ca4000(RW)
  0x1c9: frame@f9ca3000(RW)
  0x1ca: frame@f9ca2000(RW)
  0x1cb: frame@f9ca1000(RW)
  0x1cc: frame@f9ca0000(RW)
  0x1cd: frame@f9c9f000(RW)
  0x1ce: frame@f9c9e000(RW)
  0x1cf: frame@f9c9d000(RW)
  0x1d0: frame@f9c9c000(RW)
  0x1d1: frame@f9c9b000(RW)
  0x1d2: frame@f9c9a000(RW)
  0x1d3: frame@f9c99000(RW)
  0x1d4: frame@f9c98000(RW)
  0x1d5: frame@f9c97000(RW)
  0x1d6: frame@f9c96000(RW)
  0x1d7: frame@f9c95000(RW)
  0x1d8: frame@f9c94000(RW)
  0x1d9: frame@f9c93000(RW)
  0x1da: frame@f9c92000(RW)
  0x1db: frame@f9c91000(RW)
  0x1dc: frame@f9c90000(RW)
  0x1dd: frame@f9c8f000(RW)
  0x1de: frame@f9c8e000(RW)
  0x1df: frame@f9c8d000(RW)
  0x1e0: frame@f9c8c000(RW)
  0x1e1: frame@f9c8b000(RW)
  0x1e2: frame@f9c8a000(RW)
  0x1e3: frame@f9c89000(RW)
  0x1e4: frame@f9c88000(RW)
  0x1e5: frame@f9c87000(RW)
  0x1e6: frame@f9c86000(RW)
  0x1e7: frame@f9c85000(RW)
  0x1e8: frame@f9c84000(RW)
  0x1e9: frame@f9c83000(RW)
  0x1ea: frame@f9c82000(RW)
  0x1eb: frame@f9c81000(RW)
  0x1ec: frame@f9c80000(RW)
  0x1ed: frame@f9c7f000(RW)
  0x1ee: frame@f9c7e000(RW)
  0x1ef: frame@f9c7d000(RW)
  0x1f0: frame@f9c7c000(RW)
  0x1f1: frame@f9c7b000(RW)
  0x1f2: frame@f9c7a000(RW)
  0x1f3: frame@f9c79000(RW)
  0x1f4: frame@f9c78000(RW)
  0x1f5: frame@f9c77000(RW)
  0x1f6: frame@f9c76000(RW)
  0x1f7: frame@f9c75000(RW)
  0x1f8: frame@f9c74000(RW)
  0x1f9: frame@f9c73000(RW)
  0x1fa: frame@f9c72000(RW)
  0x1fb: frame@f9c71000(RW)
  0x1fc: frame@f9c70000(RW)
  0x1fd: frame@f9c6f000(RW)
  0x1fe: frame@f9c6e000(RW)
  0x1ff: frame@f9c6d000(RW)
  0x200: frame@f9c6c000(RW)
  0x201: frame@f9c6b000(RW)
  0x202: frame@f9c6a000(RW)
  0x203: frame@f9c69000(RW)
  0x204: frame@f9c68000(RW)
  0x205: frame@f9c67000(RW)
  0x206: frame@f9c66000(RW)
  0x207: frame@f9c65000(RW)
  0x208: frame@f9c64000(RW)
  0x209: frame@f9c63000(RW)
  0x20a: frame@f9c62000(RW)
  0x20b: frame@f9c61000(RW)
  0x20c: frame@f9c60000(RW)
  0x20d: frame@f9c5f000(RW)
  0x20e: frame@f9c5e000(RW)
  0x20f: frame@f9c5d000(RW)
  0x210: frame@f9c5c000(RW)
  0x211: frame@f9c5b000(RW)
  0x212: frame@f9c5a000(RW)
  0x213: frame@f9c59000(RW)
  0x214: frame@f9c58000(RW)
  0x215: frame@f9c57000(RW)
  0x216: frame@f9c56000(RW)
  0x217: frame@f9c55000(RW)
  0x218: frame@f9c54000(RW)
  0x219: frame@f9c53000(RW)
  0x21a: frame@f9c52000(RW)
  0x21b: frame@f9c51000(RW)
  0x21c: frame@f9c50000(RW)
  0x21d: frame@f9c4f000(RW)
  0x21e: frame@f9c4e000(RW)
  0x21f: frame@f9c4d000(RW)
  0x220: frame@f9c4c000(RW)
  0x221: frame@f9c4b000(RW)
  0x222: frame@f9c4a000(RW)
  0x223: frame@f9c49000(RW)
  0x224: frame@f9c48000(RW)
  0x225: frame@f9c47000(RW)
  0x226: frame@f9c46000(RW)
  0x227: frame@f9c45000(RW)
  0x228: frame@f9c44000(RW)
  0x229: frame@f9c43000(RW)
  0x22a: frame@f9c42000(RW)
  0x22b: frame@f9c41000(RW)
  0x22c: frame@f9c40000(RW)
  0x22d: frame@f9c3f000(RW)
  0x22e: frame@f9c3e000(RW)
  0x22f: frame@f9c3d000(RW)
  0x230: frame@f9c3c000(RW)
  0x231: frame@f9c3b000(RW)
  0x232: frame@f9c3a000(RW)
  0x233: frame@f9c39000(RW)
  0x234: frame@f9c38000(RW)
  0x235: frame@f9c37000(RW)
  0x236: frame@f9c36000(RW)
  0x237: frame@f9c35000(RW)
  0x238: frame@f9c34000(RW)
  0x239: frame@f9c33000(RW)
  0x23a: frame@f9c32000(RW)
  0x23b: frame@f9c31000(RW)
  0x23c: frame@f9c30000(RW)
  0x23d: frame@f9c2f000(RW)
  0x23e: frame@f9c2e000(RW)
  0x23f: frame@f9c2d000(RW)
  0x240: frame@f9c2c000(RW)
  0x241: frame@f9c2b000(RW)
  0x242: frame@f9c2a000(RW)
  0x243: frame@f9c29000(RW)
  0x244: frame@f9c28000(RW)
  0x245: frame@f9c27000(RW)
  0x246: frame@f9c26000(RW)
  0x247: frame@f9c25000(RW)
  0x248: frame@f9c24000(RW)
  0x249: frame@f9c23000(RW)
  0x24a: frame@f9c22000(RW)
  0x24b: frame@f9c21000(RW)
  0x24c: frame@f9c20000(RW)
  0x24d: frame@f9c1f000(RW)
  0x24e: frame@f9c1e000(RW)
  0x24f: frame@f9c1d000(RW)
  0x250: frame@f9c1c000(RW)
  0x251: frame@f9c1b000(RW)
  0x252: frame@f9c1a000(RW)
  0x253: frame@f9c19000(RW)
  0x254: frame@f9c18000(RW)
  0x255: frame@f9c17000(RW)
  0x256: frame@f9c16000(RW)
  0x257: frame@f9c15000(RW)
  0x258: frame@f9c14000(RW)
  0x259: frame@f9c13000(RW)
  0x25a: frame@f9c12000(RW)
  0x25b: frame@f9c11000(RW)
  0x25c: frame@f9c10000(RW)
  0x25d: frame@f9c0f000(RW)
  0x25e: frame@f9c0e000(RW)
  0x25f: frame@f9c0d000(RW)
  0x260: frame@f9c0c000(RW)
  0x261: frame@f9c0b000(RW)
  0x262: frame@f9c0a000(RW)
  0x263: frame@f9c09000(RW)
  0x264: frame@f9c08000(RW)
  0x265: frame@f9c07000(RW)
  0x266: frame@f9c06000(RW)
  0x267: frame@f9c05000(RW)
  0x268: frame@f9c04000(RW)
  0x269: frame@f9c03000(RW)
  0x26a: frame@f9c02000(RW)
  0x26b: frame@f9c01000(RW)
  0x26c: frame@f9c00000(RW)
  0x26d: frame@f9dff000(RW)
  0x26e: frame@f9dfe000(RW)
  0x26f: frame@f9dfd000(RW)
  0x270: frame@f9dfc000(RW)
  0x271: frame@f9dfb000(RW)
  0x272: frame@f9dfa000(RW)
  0x273: frame@f9df9000(RW)
  0x274: frame@f9df8000(RW)
  0x275: frame@f9df7000(RW)
  0x276: frame@f9df6000(RW)
  0x277: frame@f9df5000(RW)
  0x278: frame@f9df4000(RW)
  0x279: frame@f9df3000(RW)
  0x27a: frame@f9df2000(RW)
  0x27b: frame@f9df1000(RW)
  0x27c: frame@f9df0000(RW)
  0x27d: frame@f9def000(RW)
  0x27e: frame@f9dee000(RW)
  0x27f: frame@f9ded000(RW)
  0x280: frame@f9dec000(RW)
  0x281: frame@f9deb000(RW)
  0x282: frame@f9dea000(RW)
  0x283: frame@f9de9000(RW)
  0x284: frame@f9de8000(RW)
  0x285: frame@f9de7000(RW)
  0x286: frame@f9de6000(RW)
  0x287: frame@f9de5000(RW)
  0x288: frame@f9de4000(RW)
  0x289: frame@f9de3000(RW)
  0x28a: frame@f9de2000(RW)
  0x28b: frame@f9de1000(RW)
  0x28c: frame@f9de0000(RW)
  0x28d: frame@f9ddf000(RW)
  0x28e: frame@f9dde000(RW)
  0x28f: frame@f9ddd000(RW)
  0x290: frame@f9ddc000(RW)
  0x291: frame@f9ddb000(RW)
  0x292: frame@f9dda000(RW)
  0x293: frame@f9dd9000(RW)
  0x294: frame@f9dd8000(RW)
  0x295: frame@f9dd7000(RW)
  0x296: frame@f9dd6000(RW)
  0x297: frame@f9dd5000(RW)
  0x298: frame@f9dd4000(RW)
  0x299: frame@f9dd3000(RW)
  0x29a: frame@f9dd2000(RW)
  0x29b: frame@f9dd1000(RW)
  0x29c: frame@f9dd0000(RW)
  0x29d: frame@f9dcf000(RW)
  0x29e: frame@f9dce000(RW)
  0x29f: frame@f9dcd000(RW)
  0x2a0: frame@f9dcc000(RW)
  0x2a1: frame@f9dcb000(RW)
  0x2a2: frame@f9dca000(RW)
  0x2a3: frame@f9dc9000(RW)
}
pt@f6df8000{
  0xd0: frame@f729c000(R )
  0xd1: frame@f729b000(R )
  0xd2: frame@f729a000(R )
  0xd3: frame@f7299000(R )
  0xd4: frame@f7298000(R )
  0xd5: frame@f7297000(R )
  0xd6: frame@f7296000(R )
  0xd7: frame@f7295000(R )
  0xd8: frame@f7294000(R )
  0xd9: frame@f7293000(R )
  0xda: frame@f7292000(R )
  0xdb: frame@f7291000(R )
  0xdc: frame@f7290000(R )
  0xdd: frame@f728f000(R )
  0xde: frame@f728e000(R )
  0xdf: frame@f728d000(R )
  0xe0: frame@f728c000(R )
  0xe1: frame@f728b000(R )
  0xe2: frame@f728a000(R )
  0xe3: frame@f7289000(R )
  0xe4: frame@f7288000(R )
  0xe5: frame@f7287000(R )
  0xe6: frame@f7286000(R )
  0xe7: frame@f7285000(R )
  0xe8: frame@f7284000(R )
  0xe9: frame@f7283000(R )
  0xea: frame@f7282000(R )
  0xeb: frame@f7281000(R )
  0xec: frame@f7280000(R )
  0xed: frame@f727f000(R )
  0xee: frame@f727e000(R )
  0xef: frame@f727d000(R )
  0xf0: frame@f727c000(R )
  0xf1: frame@f727b000(R )
  0xf2: frame@f727a000(R )
  0xf3: frame@f7279000(R )
  0xf4: frame@f7278000(R )
  0xf5: frame@f7277000(R )
  0xf6: frame@f7276000(R )
  0xf7: frame@f7275000(R )
  0xf8: frame@f7274000(R )
  0xf9: frame@f7273000(R )
  0xfa: frame@f7272000(R )
  0xfb: frame@f7271000(R )
  0xfc: frame@f7270000(R )
  0xfd: frame@f726f000(R )
  0xfe: frame@f726e000(R )
  0xff: frame@f726d000(R )
  0x100: frame@f726c000(R )
  0x101: frame@f726b000(R )
  0x102: frame@f726a000(R )
  0x103: frame@f7269000(R )
  0x104: frame@f7268000(R )
  0x105: frame@f7267000(R )
  0x106: frame@f7266000(R )
  0x107: frame@f7265000(R )
  0x108: frame@f7264000(R )
  0x109: frame@f7263000(R )
  0x10a: frame@f7262000(R )
  0x10b: frame@f7261000(R )
  0x10c: frame@f7260000(R )
  0x10d: frame@f725f000(R )
  0x10e: frame@f725e000(R )
  0x10f: frame@f725d000(R )
  0x110: frame@f725c000(R )
  0x111: frame@f725b000(R )
  0x112: frame@f725a000(R )
  0x113: frame@f7259000(R )
  0x114: frame@f7258000(R )
  0x115: frame@f7257000(R )
  0x116: frame@f7256000(R )
  0x117: frame@f7255000(R )
  0x118: frame@f7254000(R )
  0x119: frame@f7253000(R )
  0x11a: frame@f7252000(R )
  0x11b: frame@f7251000(R )
  0x11c: frame@f7250000(R )
  0x11d: frame@f724f000(R )
  0x11e: frame@f724e000(R )
  0x11f: frame@f724d000(R )
  0x120: frame@f724c000(R )
  0x121: frame@f724b000(R )
  0x122: frame@f724a000(R )
  0x123: frame@f7249000(R )
  0x124: frame@f7248000(R )
  0x125: frame@f7247000(R )
  0x126: frame@f7246000(R )
  0x127: frame@f7245000(R )
  0x128: frame@f7244000(R )
  0x129: frame@f7243000(R )
  0x12a: frame@f7242000(R )
  0x12b: frame@f7241000(R )
  0x12c: frame@f7240000(R )
  0x12d: frame@f723f000(R )
  0x12e: frame@f723e000(R )
  0x12f: frame@f723d000(R )
  0x130: frame@f723c000(R )
  0x131: frame@f723b000(R )
  0x132: frame@f723a000(R )
  0x133: frame@f7239000(R )
  0x134: frame@f7238000(R )
  0x135: frame@f7237000(R )
  0x136: frame@f7236000(R )
  0x137: frame@f7235000(R )
  0x138: frame@f7234000(R )
  0x139: frame@f7233000(R )
  0x13a: frame@f7232000(R )
  0x13b: frame@f7231000(R )
  0x13c: frame@f7230000(R )
  0x13d: frame@f722f000(R )
  0x13e: frame@f722e000(R )
  0x13f: frame@f722d000(R )
  0x140: frame@f722c000(R )
  0x141: frame@f722b000(R )
  0x142: frame@f722a000(R )
  0x143: frame@f7229000(R )
  0x144: frame@f7228000(R )
  0x145: frame@f7227000(R )
  0x146: frame@f7226000(R )
  0x147: frame@f7225000(R )
  0x148: frame@f7224000(R )
  0x149: frame@f7223000(R )
  0x14a: frame@f7222000(R )
  0x14b: frame@f7221000(R )
  0x14c: frame@f7220000(R )
  0x14d: frame@f721f000(R )
  0x14e: frame@f721e000(R )
  0x14f: frame@f721d000(R )
  0x150: frame@f721c000(R )
  0x151: frame@f721b000(R )
  0x152: frame@f721a000(R )
  0x153: frame@f7219000(R )
  0x154: frame@f7218000(R )
  0x155: frame@f7217000(R )
  0x156: frame@f7216000(R )
  0x157: frame@f7215000(R )
  0x158: frame@f7214000(R )
  0x159: frame@f7213000(R )
  0x15a: frame@f7212000(R )
  0x15b: frame@f7211000(R )
  0x15c: frame@f7210000(R )
  0x15d: frame@f720f000(R )
  0x15e: frame@f720e000(R )
  0x15f: frame@f720d000(R )
  0x160: frame@f720c000(R )
  0x161: frame@f720b000(R )
  0x162: frame@f720a000(R )
  0x163: frame@f7209000(R )
  0x164: frame@f7208000(R )
  0x165: frame@f7207000(R )
  0x166: frame@f7206000(R )
  0x167: frame@f7205000(R )
  0x168: frame@f7204000(R )
  0x169: frame@f7203000(R )
  0x16a: frame@f7202000(R )
  0x16b: frame@f7201000(R )
  0x16c: frame@f7200000(R )
  0x16d: frame@f98ff000(R )
  0x16e: frame@f98fe000(R )
  0x16f: frame@f98fd000(R )
  0x170: frame@f98fc000(R )
  0x171: frame@f98fb000(R )
  0x172: frame@f98fa000(R )
  0x173: frame@f98f9000(R )
  0x174: frame@f98f8000(R )
  0x175: frame@f98f7000(R )
  0x176: frame@f98f6000(R )
  0x177: frame@f98f5000(R )
  0x178: frame@f98f4000(R )
  0x179: frame@f98f3000(R )
  0x17a: frame@f98f2000(R )
  0x17b: frame@f98f1000(R )
  0x17c: frame@f98f0000(R )
  0x17d: frame@f98ef000(R )
  0x17e: frame@f98ee000(R )
  0x17f: frame@f98ed000(R )
  0x180: frame@f98ec000(R )
  0x181: frame@f98eb000(R )
  0x182: frame@f98ea000(R )
  0x183: frame@f98e9000(R )
  0x184: frame@f98e8000(R )
  0x185: frame@f98e7000(R )
  0x186: frame@f98e6000(R )
  0x187: frame@f98e5000(R )
  0x188: frame@f98e4000(R )
  0x189: frame@f98e3000(R )
  0x18a: frame@f98e2000(R )
  0x18b: frame@f98e1000(R )
  0x18c: frame@f98e0000(R )
  0x18d: frame@f98df000(R )
  0x18e: frame@f98de000(R )
  0x18f: frame@f98dd000(R )
  0x190: frame@f98dc000(R )
  0x191: frame@f98db000(R )
  0x192: frame@f98da000(R )
  0x193: frame@f98d9000(R )
  0x194: frame@f98d8000(R )
  0x195: frame@f98d7000(R )
  0x196: frame@f98d6000(R )
  0x197: frame@f98d5000(R )
  0x198: frame@f98d4000(R )
  0x199: frame@f98d3000(R )
  0x19a: frame@f98d2000(R )
  0x19b: frame@f98d1000(R )
  0x19c: frame@f98d0000(R )
  0x19d: frame@f98cf000(R )
  0x19e: frame@f98ce000(R )
  0x19f: frame@f98cd000(R )
  0x1a0: frame@f98cc000(R )
  0x1a1: frame@f98cb000(R )
  0x1a2: frame@f98ca000(R )
  0x1a3: frame@f98c9000(R )
  0x1a4: frame@f98c8000(R )
  0x1a5: frame@f98c7000(R )
  0x1a6: frame@f98c6000(R )
  0x1a7: frame@f98c5000(R )
  0x1a8: frame@f98c4000(R )
  0x1a9: frame@f98c3000(R )
  0x1aa: frame@f98c2000(R )
  0x1ab: frame@f98c1000(R )
  0x1ac: frame@f98c0000(R )
  0x1ad: frame@f98bf000(R )
  0x1ae: frame@f98be000(R )
  0x1af: frame@f98bd000(R )
  0x1b0: frame@f98bc000(R )
  0x1b1: frame@f98bb000(R )
  0x1b2: frame@f98ba000(R )
  0x1b3: frame@f98b9000(R )
  0x1b4: frame@f98b8000(R )
  0x1b5: frame@f98b7000(R )
  0x1b6: frame@f98b6000(R )
  0x1b7: frame@f98b5000(R )
  0x1b8: frame@f98b4000(R )
  0x1b9: frame@f98b3000(R )
  0x1ba: frame@f98b2000(R )
  0x1bb: frame@f98b1000(R )
  0x1bc: frame@f98b0000(R )
  0x1bd: frame@f98af000(R )
  0x1be: frame@f98ae000(R )
  0x1bf: frame@f98ad000(R )
  0x1c0: frame@f98ac000(R )
  0x1c1: frame@f98ab000(R )
  0x1c2: frame@f98aa000(R )
  0x1c3: frame@f98a9000(R )
  0x1c4: frame@f98a8000(R )
  0x1c5: frame@f98a7000(R )
  0x1c6: frame@f98a6000(R )
  0x1c7: frame@f98a5000(R )
  0x1c8: frame@f98a4000(R )
  0x1c9: frame@f98a3000(R )
  0x1ca: frame@f98a2000(R )
  0x1cb: frame@f98a1000(R )
  0x1cc: frame@f98a0000(R )
  0x1cd: frame@f989f000(R )
  0x1ce: frame@f989e000(R )
  0x1cf: frame@f989d000(R )
  0x1d0: frame@f989c000(R )
  0x1d1: frame@f989b000(R )
  0x1d2: frame@f989a000(R )
  0x1d3: frame@f9899000(R )
  0x1d4: frame@f9898000(R )
  0x1d5: frame@f9897000(R )
  0x1d6: frame@f9896000(R )
  0x1d7: frame@f9895000(R )
  0x1d8: frame@f9894000(R )
  0x1d9: frame@f9893000(R )
  0x1da: frame@f9892000(R )
  0x1db: frame@f9891000(R )
  0x1dc: frame@f9890000(R )
  0x1dd: frame@f988f000(R )
  0x1de: frame@f988e000(R )
  0x1df: frame@f988d000(R )
  0x1e0: frame@f988c000(R )
  0x1e1: frame@f988b000(R )
  0x1e2: frame@f988a000(R )
  0x1e3: frame@f9889000(R )
  0x1e4: frame@f9888000(R )
  0x1e5: frame@f9887000(R )
  0x1e6: frame@f9886000(R )
  0x1e7: frame@f9885000(R )
  0x1e8: frame@f9884000(R )
  0x1e9: frame@f9883000(R )
  0x1ea: frame@f9882000(R )
  0x1eb: frame@f9881000(R )
  0x1ec: frame@f9880000(R )
  0x1ed: frame@f987f000(R )
  0x1ee: frame@f987e000(R )
  0x1ef: frame@f987d000(R )
  0x1f0: frame@f987c000(R )
  0x1f1: frame@f987b000(R )
  0x1f2: frame@f987a000(R )
  0x1f3: frame@f9879000(R )
  0x1f4: frame@f9878000(R )
  0x1f5: frame@f9877000(R )
  0x1f6: frame@f9876000(R )
  0x1f7: frame@f9875000(R )
  0x1f8: frame@f9874000(R )
  0x1f9: frame@f9873000(R )
  0x1fa: frame@f9872000(R )
  0x1fb: frame@f9871000(R )
  0x1fc: frame@f9870000(R )
  0x1fd: frame@f986f000(R )
  0x1fe: frame@f986e000(R )
  0x1ff: frame@f986d000(R )
  0x200: frame@f986c000(R )
  0x201: frame@f986b000(R )
  0x202: frame@f986a000(R )
  0x203: frame@f9869000(R )
  0x204: frame@f9868000(R )
  0x205: frame@f9867000(R )
  0x206: frame@f9866000(R )
  0x207: frame@f9865000(R )
  0x208: frame@f9864000(R )
  0x209: frame@f9863000(R )
  0x20a: frame@f9862000(R )
  0x20b: frame@f9861000(R )
  0x20c: frame@f9860000(R )
  0x20d: frame@f985f000(R )
  0x20e: frame@f985e000(R )
  0x20f: frame@f985d000(R )
  0x210: frame@f985c000(R )
  0x211: frame@f985b000(R )
  0x212: frame@f985a000(R )
  0x213: frame@f9859000(R )
  0x214: frame@f9858000(R )
  0x215: frame@f9857000(R )
  0x216: frame@f9856000(R )
  0x217: frame@f9855000(R )
  0x218: frame@f9854000(R )
  0x219: frame@f9853000(R )
  0x21a: frame@f9852000(R )
  0x21b: frame@f9851000(R )
  0x21c: frame@f9850000(R )
  0x21d: frame@f984f000(R )
  0x21e: frame@f984e000(R )
  0x21f: frame@f984d000(R )
  0x220: frame@f984c000(R )
  0x221: frame@f984b000(R )
  0x222: frame@f984a000(R )
  0x223: frame@f9849000(R )
  0x224: frame@f9848000(R )
  0x225: frame@f9847000(R )
  0x226: frame@f9846000(R )
  0x227: frame@f9845000(R )
  0x228: frame@f9844000(R )
  0x229: frame@f9843000(R )
  0x22a: frame@f9842000(R )
  0x22b: frame@f9841000(R )
  0x22c: frame@f9840000(R )
  0x22d: frame@f983f000(R )
  0x22e: frame@f983e000(R )
  0x22f: frame@f983d000(R )
  0x230: frame@f983c000(R )
  0x231: frame@f983b000(R )
  0x232: frame@f983a000(R )
  0x233: frame@f9839000(R )
  0x234: frame@f9838000(R )
  0x235: frame@f9837000(R )
  0x236: frame@f9836000(R )
  0x237: frame@f9835000(R )
  0x238: frame@f9834000(R )
  0x239: frame@f9833000(R )
  0x23a: frame@f9832000(R )
  0x23b: frame@f9831000(R )
  0x23c: frame@f9830000(R )
  0x23d: frame@f982f000(R )
  0x23e: frame@f982e000(R )
  0x23f: frame@f982d000(R )
  0x240: frame@f982c000(R )
  0x241: frame@f982b000(R )
  0x242: frame@f982a000(R )
  0x243: frame@f9829000(R )
  0x244: frame@f9828000(R )
  0x245: frame@f9827000(R )
  0x246: frame@f9826000(R )
  0x247: frame@f9825000(R )
  0x248: frame@f9824000(R )
  0x249: frame@f9823000(R )
  0x24a: frame@f9822000(R )
  0x24b: frame@f9821000(R )
  0x24c: frame@f9820000(R )
  0x24d: frame@f981f000(R )
  0x24e: frame@f981e000(R )
  0x24f: frame@f981d000(R )
  0x250: frame@f981c000(R )
  0x251: frame@f981b000(R )
  0x252: frame@f981a000(R )
  0x253: frame@f9819000(R )
  0x254: frame@f9818000(R )
  0x255: frame@f9817000(R )
  0x256: frame@f9816000(R )
  0x257: frame@f9815000(R )
  0x258: frame@f9814000(R )
  0x259: frame@f9813000(R )
  0x25a: frame@f9812000(R )
  0x25b: frame@f9811000(R )
  0x25c: frame@f9810000(R )
  0x25d: frame@f980f000(R )
  0x25e: frame@f980e000(R )
  0x25f: frame@f980d000(R )
  0x260: frame@f980c000(R )
  0x261: frame@f980b000(R )
  0x262: frame@f980a000(R )
  0x263: frame@f9809000(R )
  0x264: frame@f9808000(R )
  0x265: frame@f9807000(R )
  0x266: frame@f9806000(R )
  0x267: frame@f9805000(R )
  0x268: frame@f9804000(R )
  0x269: frame@f9803000(R )
  0x26a: frame@f9802000(R )
  0x26b: frame@f9801000(R )
  0x26c: frame@f9800000(R )
  0x26d: frame@f99ff000(R )
  0x26e: frame@f99fe000(R )
  0x26f: frame@f99fd000(R )
  0x270: frame@f99fc000(R )
  0x271: frame@f99fb000(R )
  0x272: frame@f99fa000(R )
  0x273: frame@f99f9000(R )
  0x274: frame@f99f8000(R )
  0x275: frame@f99f7000(R )
  0x276: frame@f99f6000(R )
  0x277: frame@f99f5000(R )
  0x278: frame@f99f4000(R )
  0x279: frame@f99f3000(R )
  0x27a: frame@f99f2000(R )
  0x27b: frame@f99f1000(R )
  0x27c: frame@f99f0000(R )
  0x27d: frame@f99ef000(R )
  0x27e: frame@f99ee000(R )
  0x27f: frame@f99ed000(R )
  0x280: frame@f99ec000(R )
  0x281: frame@f99eb000(R )
  0x282: frame@f99ea000(R )
  0x283: frame@f99e9000(R )
  0x284: frame@f99e8000(R )
  0x285: frame@f99e7000(R )
  0x286: frame@f99e6000(R )
  0x287: frame@f99e5000(R )
  0x288: frame@f99e4000(R )
  0x289: frame@f99e3000(R )
  0x28a: frame@f99e2000(R )
  0x28b: frame@f99e1000(R )
  0x28c: frame@f99e0000(R )
  0x28d: frame@f99df000(R )
  0x28e: frame@f99de000(R )
  0x28f: frame@f99dd000(R )
  0x290: frame@f99dc000(R )
  0x291: frame@f99db000(R )
  0x292: frame@f99da000(R )
  0x293: frame@f99d9000(R )
  0x294: frame@f99d8000(R )
  0x295: frame@f99d7000(R )
  0x296: frame@f99d6000(R )
  0x297: frame@f99d5000(R )
  0x298: frame@f99d4000(R )
  0x299: frame@f99d3000(R )
  0x29a: frame@f99d2000(R )
  0x29b: frame@f99d1000(R )
  0x29c: frame@f99d0000(R )
  0x29d: frame@f99cf000(R )
  0x29e: frame@f99ce000(R )
  0x29f: frame@f99cd000(R )
  0x2a0: frame@f99cc000(R )
  0x2a1: frame@f99cb000(R )
  0x2a2: frame@f99ca000(R )
  0x2a3: frame@f99c9000(R )
  0x2a4: frame@f99c8000(R )
  0x2a5: frame@f99c7000(R )
  0x2a6: frame@f99c6000(R )
  0x2a7: frame@f99c5000(R )
  0x2a8: frame@f99c4000(R )
  0x2a9: frame@f99c3000(R )
  0x2aa: frame@f99c2000(R )
  0x2ab: frame@f99c1000(R )
  0x2ac: frame@f99c0000(R )
  0x2ad: frame@f99bf000(R )
  0x2ae: frame@f99be000(R )
  0x2af: frame@f99bd000(R )
  0x2b0: frame@f99bc000(R )
  0x2b1: frame@f99bb000(R )
  0x2b2: frame@f99ba000(R )
  0x2b3: frame@f99b9000(R )
  0x2b4: frame@f99b8000(R )
  0x2b5: frame@f99b7000(R )
  0x2b6: frame@f99b6000(R )
  0x2b7: frame@f99b5000(R )
  0x2b8: frame@f99b4000(R )
  0x2b9: frame@f99b3000(R )
  0x2ba: frame@f99b2000(R )
  0x2bb: frame@f99b1000(R )
  0x2bc: frame@f99b0000(R )
  0x2bd: frame@f99af000(R )
  0x2be: frame@f99ae000(R )
  0x2bf: frame@f99ad000(R )
  0x2c0: frame@f99ac000(R )
  0x2c1: frame@f99ab000(R )
  0x2c2: frame@f99aa000(R )
  0x2c3: frame@f99a9000(R )
  0x2c4: frame@f99a8000(R )
  0x2c5: frame@f99a7000(R )
  0x2c6: frame@f99a6000(R )
  0x2c7: frame@f99a5000(R )
  0x2c8: frame@f99a4000(R )
  0x2c9: frame@f99a3000(R )
  0x2ca: frame@f99a2000(R )
  0x2cb: frame@f99a1000(R )
  0x2cc: frame@f99a0000(R )
  0x2cd: frame@f999f000(R )
  0x2ce: frame@f999e000(R )
  0x2cf: frame@f999d000(R )
  0x2d0: frame@f999c000(R )
  0x2d1: frame@f999b000(R )
  0x2d2: frame@f999a000(R )
  0x2d3: frame@f9999000(R )
  0x2d4: frame@f9998000(R )
  0x2d5: frame@f9997000(R )
  0x2d6: frame@f9996000(R )
  0x2d7: frame@f9995000(R )
  0x2d8: frame@f9994000(R )
  0x2d9: frame@f9993000(R )
  0x2da: frame@f9992000(R )
  0x2db: frame@f9991000(R )
  0x2dc: frame@f9990000(R )
  0x2dd: frame@f998f000(R )
  0x2de: frame@f998e000(R )
  0x2df: frame@f998d000(R )
  0x2e0: frame@f998c000(R )
  0x2e1: frame@f998b000(R )
  0x2e2: frame@f998a000(R )
  0x2e3: frame@f9989000(R )
  0x2e4: frame@f9988000(R )
  0x2e5: frame@f9987000(R )
  0x2e6: frame@f9986000(R )
  0x2e7: frame@f9985000(R )
  0x2e8: frame@f9984000(R )
  0x2e9: frame@f9983000(R )
  0x2ea: frame@f9982000(R )
  0x2eb: frame@f9981000(R )
  0x2ec: frame@f9980000(R )
  0x2ed: frame@f997f000(R )
  0x2ee: frame@f997e000(R )
  0x2ef: frame@f997d000(R )
  0x2f0: frame@f997c000(R )
  0x2f1: frame@f997b000(R )
  0x2f2: frame@f997a000(R )
  0x2f3: frame@f9979000(R )
  0x2f4: frame@f9978000(R )
  0x2f5: frame@f9977000(R )
  0x2f6: frame@f9976000(RW)
  0x2f7: frame@f9975000(RW)
  0x2f8: frame@f9974000(RW)
  0x2f9: frame@f9973000(RW)
  0x2fa: frame@f9972000(RW)
  0x2fb: frame@f9971000(RW)
  0x2fc: frame@f9970000(RW)
  0x2fd: frame@f996f000(RW)
  0x2fe: frame@f996e000(RW)
  0x2ff: frame@f996d000(RW)
  0x300: frame@f996c000(RW)
  0x301: frame@f996b000(RW)
  0x302: frame@f996a000(RW)
  0x303: frame@f9969000(RW)
  0x304: frame@f9968000(RW)
  0x305: frame@f9967000(RW)
  0x306: frame@f9966000(RW)
  0x307: frame@f9965000(RW)
  0x308: frame@f9964000(RW)
  0x309: frame@f9963000(RW)
  0x30a: frame@f9962000(RW)
  0x30b: frame@f9961000(RW)
  0x30c: frame@f9960000(RW)
  0x30d: frame@f995f000(RW)
  0x30e: frame@f995e000(RW)
  0x30f: frame@f995d000(RW)
  0x310: frame@f995c000(RW)
  0x311: frame@f995b000(RW)
  0x312: frame@f995a000(RW)
  0x313: frame@f9959000(RW)
  0x314: frame@f9958000(RW)
  0x315: frame@f9957000(RW)
  0x316: frame@f9956000(RW)
  0x317: frame@f9955000(RW)
  0x318: frame@f9954000(RW)
  0x319: frame@f9953000(RW)
  0x31a: frame@f9952000(RW)
  0x31b: frame@f9951000(RW)
  0x31c: frame@f9950000(RW)
  0x31d: frame@f994f000(RW)
  0x31e: frame@f994e000(RW)
  0x31f: frame@f994d000(RW)
  0x320: frame@f994c000(RW)
  0x321: frame@f994b000(RW)
  0x322: frame@f994a000(RW)
  0x323: frame@f9949000(RW)
  0x324: frame@f9948000(RW)
  0x325: frame@f9947000(RW)
  0x326: frame@f9946000(RW)
  0x327: frame@f9945000(RW)
  0x328: frame@f9944000(RW)
  0x329: frame@f9943000(RW)
  0x32a: frame@f9942000(RW)
  0x32b: frame@f9941000(RW)
  0x32c: frame@f9940000(RW)
  0x32d: frame@f993f000(RW)
  0x32e: frame@f993e000(RW)
  0x32f: frame@f993d000(RW)
  0x330: frame@f993c000(RW)
  0x331: frame@f993b000(RW)
  0x332: frame@f993a000(RW)
  0x333: frame@f9939000(RW)
  0x334: frame@f9938000(RW)
  0x335: frame@f9937000(RW)
  0x336: frame@f9936000(RW)
  0x337: frame@f9935000(RW)
  0x338: frame@f9934000(RW)
  0x339: frame@f9933000(RW)
  0x33a: frame@f9932000(RW)
  0x33b: frame@f9931000(RW)
  0x33c: frame@f9930000(RW)
  0x33d: frame@f992f000(RW)
  0x33e: frame@f992e000(RW)
  0x33f: frame@f992d000(RW)
  0x340: frame@f992c000(RW)
  0x341: frame@f992b000(RW)
  0x342: frame@f992a000(RW)
  0x343: frame@f9929000(RW)
  0x344: frame@f9928000(RW)
  0x345: frame@f9927000(RW)
  0x346: frame@f9926000(RW)
  0x347: frame@f9925000(RW)
  0x348: frame@f9924000(RW)
  0x349: frame@f9923000(RW)
  0x34a: frame@f9922000(RW)
  0x34b: frame@f9921000(RW)
  0x34c: frame@f9920000(RW)
  0x34d: frame@f991f000(RW)
  0x34e: frame@f991e000(RW)
  0x34f: frame@f991d000(RW)
  0x350: frame@f991c000(RW)
  0x351: frame@f991b000(RW)
  0x352: frame@f991a000(RW)
  0x353: frame@f9919000(RW)
  0x354: frame@f9918000(RW)
  0x355: frame@f9917000(RW)
  0x356: frame@f9916000(RW)
  0x357: frame@f9915000(RW)
  0x358: frame@f9914000(RW)
  0x359: frame@f9913000(RW)
  0x35a: frame@f9912000(RW)
  0x35b: frame@f9911000(RW)
  0x35c: frame@f9910000(RW)
  0x35d: frame@f990f000(RW)
  0x35e: frame@f990e000(RW)
  0x35f: frame@f990d000(RW)
  0x360: frame@f990c000(RW)
  0x361: frame@f990b000(RW)
  0x362: frame@f990a000(RW)
  0x363: frame@f9909000(RW)
  0x364: frame@f9908000(RW)
  0x365: frame@f9907000(RW)
  0x366: frame@f9906000(RW)
  0x367: frame@f9905000(RW)
  0x368: frame@f9904000(RW)
  0x369: frame@f9903000(RW)
  0x36a: frame@f9902000(RW)
  0x36b: frame@f9901000(RW)
  0x36c: frame@f9900000(RW)
  0x36d: frame@f9aff000(RW)
  0x36e: frame@f9afe000(RW)
  0x36f: frame@f9afd000(RW)
  0x370: frame@f9afc000(RW)
  0x371: frame@f9afb000(RW)
  0x372: frame@f9afa000(RW)
  0x373: frame@f9af9000(RW)
  0x374: frame@f9af8000(RW)
  0x375: frame@f9af7000(RW)
  0x376: frame@f9af6000(RW)
  0x377: frame@f9af5000(RW)
  0x378: frame@f9af4000(RW)
  0x379: frame@f9af3000(RW)
  0x37a: frame@f9af2000(RW)
  0x37b: frame@f9af1000(RW)
  0x37c: frame@f9af0000(RW)
  0x37d: frame@f9aef000(RW)
  0x37e: frame@f9aee000(RW)
  0x37f: frame@f9aed000(RW)
  0x380: frame@f9aec000(RW)
  0x381: frame@f9aeb000(RW)
  0x382: frame@f9aea000(RW)
  0x383: frame@f9ae9000(RW)
  0x384: frame@f9ae8000(RW)
  0x385: frame@f9ae7000(RW)
  0x386: frame@f9ae6000(RW)
  0x387: frame@f9ae5000(RW)
  0x388: frame@f9ae4000(RW)
  0x389: frame@f9ae3000(RW)
  0x38a: frame@f9ae2000(RW)
  0x38b: frame@f9ae1000(RW)
  0x38c: frame@f9ae0000(RW)
  0x38d: frame@f9adf000(RW)
  0x38e: frame@f9ade000(RW)
  0x38f: frame@f9add000(RW)
  0x390: frame@f9adc000(RW)
  0x391: frame@f9adb000(RW)
  0x392: frame@f9ada000(RW)
  0x393: frame@f9ad9000(RW)
  0x394: frame@f9ad8000(RW)
  0x395: frame@f9ad7000(RW)
  0x396: frame@f9ad6000(RW)
  0x397: frame@f9ad5000(RW)
  0x398: frame@f9ad4000(RW)
  0x399: frame@f9ad3000(RW)
  0x39a: frame@f9ad2000(RW)
  0x39b: frame@f9ad1000(RW)
  0x39c: frame@f9ad0000(RW)
  0x39d: frame@f9acf000(RW)
  0x39e: frame@f9ace000(RW)
  0x39f: frame@f9acd000(RW)
  0x3a0: frame@f9acc000(RW)
  0x3a1: frame@f9acb000(RW)
  0x3a2: frame@f9aca000(RW)
  0x3a3: frame@f9ac9000(RW)
  0x3a4: frame@f9ac8000(RW)
  0x3a5: frame@f9ac7000(RW)
  0x3a6: frame@f9ac6000(RW)
  0x3a7: frame@f9ac5000(RW)
  0x3a8: frame@f9ac4000(RW)
  0x3a9: frame@f9ac3000(RW)
  0x3aa: frame@f9ac2000(RW)
  0x3ab: frame@f9ac1000(RW)
  0x3ac: frame@f9ac0000(RW)
  0x3ad: frame@f9abf000(RW)
  0x3ae: frame@f9abe000(RW)
  0x3af: frame@f9abd000(RW)
  0x3b0: frame@f9abc000(RW)
  0x3b1: frame@f9abb000(RW)
  0x3b2: frame@f9aba000(RW)
  0x3b3: frame@f9ab9000(RW)
  0x3b4: frame@f9ab8000(RW)
  0x3b5: frame@f9ab7000(RW)
  0x3b6: frame@f9ab6000(RW)
  0x3b7: frame@f9ab5000(RW)
  0x3b8: frame@f9ab4000(RW)
  0x3b9: frame@f9ab3000(RW)
  0x3ba: frame@f9ab2000(RW)
  0x3bb: frame@f9ab1000(RW)
  0x3bc: frame@f9ab0000(RW)
  0x3bd: frame@f9aaf000(RW)
  0x3be: frame@f9aae000(RW)
  0x3bf: frame@f9aad000(RW)
  0x3c0: frame@f9aac000(RW)
  0x3c1: frame@f9aab000(RW)
  0x3c2: frame@f9aaa000(RW)
  0x3c3: frame@f9aa9000(RW)
  0x3c4: frame@f9aa8000(RW)
  0x3c5: frame@f9aa7000(RW)
  0x3c6: frame@f9aa6000(RW)
  0x3c7: frame@f9aa5000(RW)
  0x3c8: frame@f9aa4000(RW)
  0x3c9: frame@f9aa3000(RW)
  0x3ca: frame@f9aa2000(RW)
  0x3cb: frame@f9aa1000(RW)
  0x3cc: frame@f9aa0000(RW)
  0x3cd: frame@f9a9f000(RW)
  0x3ce: frame@f9a9e000(RW)
  0x3cf: frame@f9a9d000(RW)
  0x3d0: frame@f9a9c000(RW)
  0x3d1: frame@f9a9b000(RW)
  0x3d2: frame@f9a9a000(RW)
  0x3d3: frame@f9a99000(RW)
  0x3d4: frame@f9a98000(RW)
  0x3d5: frame@f9a97000(RW)
  0x3d6: frame@f9a96000(RW)
  0x3d7: frame@f9a95000(RW)
  0x3d8: frame@f9a94000(RW)
  0x3d9: frame@f9a93000(RW)
  0x3da: frame@f9a92000(RW)
  0x3db: frame@f9a91000(RW)
  0x3dc: frame@f9a90000(RW)
  0x3dd: frame@f9a8f000(RW)
  0x3de: frame@f9a8e000(RW)
  0x3df: frame@f9a8d000(RW)
  0x3e0: frame@f9a8c000(RW)
  0x3e1: frame@f9a8b000(RW)
  0x3e2: frame@f9a8a000(RW)
  0x3e3: frame@f9a89000(RW)
  0x3e4: frame@f9a88000(RW)
  0x3e5: frame@f9a87000(RW)
  0x3e6: frame@f9a86000(RW)
  0x3e7: frame@f9a85000(RW)
  0x3e8: frame@f9a84000(RW)
  0x3e9: frame@f9a83000(RW)
  0x3ea: frame@f9a82000(RW)
  0x3eb: frame@f9a81000(RW)
  0x3ec: frame@f9a80000(RW)
  0x3ed: frame@f9a7f000(RW)
  0x3ee: frame@f9a7e000(RW)
  0x3ef: frame@f9a7d000(RW)
  0x3f0: frame@f9a7c000(RW)
  0x3f1: frame@f9a7b000(RW)
  0x3f2: frame@f9a7a000(RW)
  0x3f3: frame@f9a79000(RW)
  0x3f4: frame@f9a78000(RW)
  0x3f5: frame@f9a77000(RW)
  0x3f6: frame@f9a76000(RW)
  0x3f7: frame@f9a75000(RW)
  0x3f8: frame@f9a74000(RW)
  0x3f9: frame@f9a73000(RW)
  0x3fa: frame@f9a72000(RW)
  0x3fb: frame@f9a71000(RW)
  0x3fc: frame@f9a70000(RW)
  0x3fd: frame@f9a6f000(RW)
  0x3fe: frame@f9a6e000(RW)
  0x3ff: frame@f9a6d000(RW)
}
